//revision : "V1.2.2"
//date : "Dec 30 2011"
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM, INC.
//Copyright (c) 2002-2009 ARM, Inc.
//The confidential and proprietary information contained in this file
//may only be used by a person authorised under and to the extent
//permitted by a subsisting licensing agreement from ARM Limited.
//
//(C) COPYRIGHT 2004-2009 ARM Limited.
//ALL RIGHTS RESERVED
//
//This entire notice must be reproduced on all copies of this file
//and copies of this file may only be made by a person if such person
//is permitted to do so under the terms of a subsisting license
//agreement from ARM Limited or Samsung Electronics.
//
//Modification of this file is not permitted for any one and any case. 
//Samsung Electronics has no responsibility for any problem caused by unpermitted modification of this file.

`define ARM_PROP_FF_DELAY 	0.3
`define ARM_PROP_DELAY 	0.01
`define ARM_INVALID_DELAY 	100.0

`define ARM_PERIOD 	0.0
`define ARM_WIDTH 	0.0
`define ARM_SETUP_TIME 	0.0
`define ARM_HOLD_TIME 	0.0
`define ARM_RECOVERY_TIME 	0.0
`define ARM_REMOVAL_TIME 	0.0
`define ARM_WIDTH_THD 	0.0

`timescale 1ns/1ps
`celldefine
module DFFQ_X0P5M_A12TR (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf #0     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
	`ifdef PRE_NETLIST_SIM
		buf #0.1  I1 (Q, n0);
	`else
	  buf     I1 (Q, n0);
	`endif

wire ENABLE_NOT_D ;
wire ENABLE_D ;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_D == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_FF_DELAY,`ARM_PROP_FF_DELAY);

endspecify
endmodule // DFFQ_X0P5M_A12TR
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ADDF_X1M_A12TR (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X1M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X0P5M_A12TR (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X0P5M_A12TR (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21A1AI2_X0P5M_A12TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  or I1(outB, outA, B0);
  nand I3(Y, outB, C0);




specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21A1AI2_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21B_X0P5M_A12TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21B_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X0P5M_A12TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X0P5M_A12TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X0P5M_A12TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X0P5M_A12TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22BB_X0P5M_A12TR (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  and I0(outA, A0, A1);
  not I1 (outB0, B0N);
  not I2 (outB1, B1N);
  and I3 (outB, outB0, outB1);
  nor I4 (Y,outA,outB);

specify
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22BB_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X0P5M_A12TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2XB1_X0P5M_A12TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2XB1_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X0P5M_A12TR (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGENI_X1M_A12TR (CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I3 (cout, a_and_b, a_and_ci, b_and_ci);
  not I4 (CON, cout);


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGENI_X1M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CGEN_X1M_A12TR (CO, A, B, CI);
output CO;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or I4 (CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CGEN_X1M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X0P5B_A12TR (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X0P5B_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XB_X0P5M_A12TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XB_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X0P5A_A12TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X0P5A_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BB_X0P5M_A12TR (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BB_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X0P5M_A12TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XB_X0P5M_A12TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XB_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X0P5B_A12TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X0P5B_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BB_X0P5M_A12TR (Y, AN, BN, C);
output Y;
input AN, BN, C;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BB_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X0P7M_A12TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X0P7M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA1B2_X0P7M_A12TR (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;



  nor I1 (outB, B0, B1);
  nor I2 (Y, A0N, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA1B2_X0P7M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA211_X0P5M_A12TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA211_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21A1OI2_X0P7M_A12TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;


  or I0(outA, A0, A1);
  and I1(outB, outA, B0);
  nor I3(Y, outB, C0);



specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21A1OI2_X0P7M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X0P5M_A12TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X0P5M_A12TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X0P5M_A12TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X0P5M_A12TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22BB_X0P5M_A12TR (Y, A0, A1, B0N, B1N);
output Y;
input A0, A1, B0N, B1N;



  not  I0 (outB0, B0N);
  not  I1 (outB1, B1N);
  or   I2 (outB, outB0, outB1);
  or   I3 (outA, A0, A1);
  nand I4 (Y, outA, outB);


specify
if (B0N==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b0 && B1N==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0N==1'b1 && B1N==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22BB_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X0P5M_A12TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X0P5M_A12TR (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X0P5M_A12TR (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X0P5M_A12TR (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X0P5M_A12TR (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X0P5M_A12TR
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X0P5M_A12TR (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X0P5M_A12TR
`endcelldefine

//20101116 udp_dff
`ifdef FF_NO_X_OUT
module udp_dff  (out, in, clk, clr_, set_, NOTIFIER);
   output out;
   input   in, clk, clr_, set_, NOTIFIER;
   reg out;
   wire pout;

   initial out <= `ForcedX_VAL;

   always @(pout) begin
   	if(pout===1'bx)
   		out <= `ForcedX_VAL;
   	else
   		out <= pout;
   end

   _udp_dff u1 (pout,   in, clk, clr_, set_, NOTIFIER);

endmodule

primitive _udp_dff  (out, in, clk, clr_, set_, NOTIFIER);
`else
primitive udp_dff (out, in, clk, clr_, set_, NOTIFIER);
`endif
   output out;  
   input  in, clk, clr_, set_, NOTIFIER;
   reg    out;

   table

// in  clk  clr_   set_  NOT  : Qt : Qt+1
//
   0  r   ?   1   ?   : ?  :  0  ; // clock in 0
   1  r   1   ?   ?   : ?  :  1  ; // clock in 1
   1  *   1   ?   ?   : 1  :  1  ; // reduce pessimism
   0  *   ?   1   ?   : 0  :  0  ; // reduce pessimism
   ?  f   ?   ?   ?   : ?  :  -  ; // no changes on negedge clk
   *  b   ?   ?   ?   : ?  :  -  ; // no changes when in switches
   ?  ?   ?   0   ?   : ?  :  1  ; // set output
   ?  b   1   *   ?   : 1  :  1  ; // cover all transistions on set_
   1  x   1   *   ?   : 1  :  1  ; // cover all transistions on set_
   ?  ?   0   1   ?   : ?  :  0  ; // reset output
   ?  b   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
   0  x   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
   ?  ?   ?   ?   *   : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_dff


module mul_add ( clk1, clk2, reset, a, b, out );
  input [31:0] a;
  input [31:0] b;
  output [31:0] out;
  input clk1, clk2, reset;
  wire   \areg_stage1/N34 , \areg_stage1/N33 , \areg_stage1/N32 ,
         \areg_stage1/N31 , \areg_stage1/N30 , \areg_stage1/N29 ,
         \areg_stage1/N28 , \areg_stage1/N27 , \areg_stage1/N26 ,
         \areg_stage1/N25 , \areg_stage1/N24 , \areg_stage1/N23 ,
         \areg_stage1/N22 , \areg_stage1/N21 , \areg_stage1/N20 ,
         \areg_stage1/N19 , \areg_stage1/N18 , \areg_stage1/N17 ,
         \areg_stage1/N16 , \areg_stage1/N15 , \areg_stage1/N14 ,
         \areg_stage1/N13 , \areg_stage1/N12 , \areg_stage1/N11 ,
         \areg_stage1/N10 , \areg_stage1/N9 , \areg_stage1/N8 ,
         \areg_stage1/N7 , \areg_stage1/N6 , \areg_stage1/N5 ,
         \areg_stage1/N4 , \areg_stage1/N3 , \breg_stage1/N34 ,
         \breg_stage1/N33 , \breg_stage1/N32 , \breg_stage1/N31 ,
         \breg_stage1/N30 , \breg_stage1/N29 , \breg_stage1/N28 ,
         \breg_stage1/N27 , \breg_stage1/N26 , \breg_stage1/N25 ,
         \breg_stage1/N24 , \breg_stage1/N23 , \breg_stage1/N22 ,
         \breg_stage1/N21 , \breg_stage1/N20 , \breg_stage1/N19 ,
         \breg_stage1/N18 , \breg_stage1/N17 , \breg_stage1/N16 ,
         \breg_stage1/N15 , \breg_stage1/N14 , \breg_stage1/N13 ,
         \breg_stage1/N12 , \breg_stage1/N11 , \breg_stage1/N10 ,
         \breg_stage1/N9 , \breg_stage1/N8 , \breg_stage1/N7 ,
         \breg_stage1/N6 , \breg_stage1/N5 , \breg_stage1/N4 ,
         \breg_stage1/N3 , \accreg_stage2/N34 , \accreg_stage2/N33 ,
         \accreg_stage2/N32 , \accreg_stage2/N31 , \accreg_stage2/N30 ,
         \accreg_stage2/N29 , \accreg_stage2/N28 , \accreg_stage2/N27 ,
         \accreg_stage2/N26 , \accreg_stage2/N25 , \accreg_stage2/N24 ,
         \accreg_stage2/N23 , \accreg_stage2/N22 , \accreg_stage2/N21 ,
         \accreg_stage2/N20 , \accreg_stage2/N19 , \accreg_stage2/N18 ,
         \accreg_stage2/N17 , \accreg_stage2/N16 , \accreg_stage2/N15 ,
         \accreg_stage2/N14 , \accreg_stage2/N13 , \accreg_stage2/N12 ,
         \accreg_stage2/N11 , \accreg_stage2/N10 , \accreg_stage2/N9 ,
         \accreg_stage2/N8 , \accreg_stage2/N7 , \accreg_stage2/N6 ,
         \accreg_stage2/N5 , \accreg_stage2/N4 , \accreg_stage2/N3 ,
         \outreg_stage2/N34 , \outreg_stage2/N33 , \outreg_stage2/N32 ,
         \outreg_stage2/N31 , \outreg_stage2/N30 , \outreg_stage2/N29 ,
         \outreg_stage2/N28 , \outreg_stage2/N27 , \outreg_stage2/N26 ,
         \outreg_stage2/N25 , \outreg_stage2/N24 , \outreg_stage2/N23 ,
         \outreg_stage2/N22 , \outreg_stage2/N21 , \outreg_stage2/N20 ,
         \outreg_stage2/N19 , \outreg_stage2/N18 , \outreg_stage2/N17 ,
         \outreg_stage2/N16 , \outreg_stage2/N15 , \outreg_stage2/N14 ,
         \outreg_stage2/N13 , \outreg_stage2/N12 , \outreg_stage2/N11 ,
         \outreg_stage2/N10 , \outreg_stage2/N9 , \outreg_stage2/N8 ,
         \outreg_stage2/N7 , \outreg_stage2/N6 , \outreg_stage2/N5 ,
         \outreg_stage2/N4 , \outreg_stage2/N3 , n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484;
  wire   [31:0] a_s1;
  wire   [31:0] b_s1;
  wire   [31:0] acc_s2;
  wire   [31:0] in_s2;

  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[14]  ( .D(\outreg_stage2/N17 ), .CK(
        clk2), .Q(in_s2[14]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[29]  ( .D(\outreg_stage2/N32 ), .CK(
        clk2), .Q(in_s2[29]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[31]  ( .D(\areg_stage1/N34 ), .CK(clk1), 
        .Q(a_s1[31]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[14]  ( .D(\accreg_stage2/N17 ), .CK(
        clk2), .Q(acc_s2[14]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[29]  ( .D(\accreg_stage2/N32 ), .CK(
        clk2), .Q(acc_s2[29]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[29]  ( .D(\areg_stage1/N32 ), .CK(clk1), 
        .Q(a_s1[29]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[17]  ( .D(\breg_stage1/N20 ), .CK(clk1), 
        .Q(b_s1[17]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[2]  ( .D(\areg_stage1/N5 ), .CK(clk1), 
        .Q(a_s1[2]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[31]  ( .D(\accreg_stage2/N34 ), .CK(
        clk2), .Q(acc_s2[31]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[1]  ( .D(\outreg_stage2/N4 ), .CK(clk2), .Q(in_s2[1]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[2]  ( .D(\outreg_stage2/N5 ), .CK(clk2), .Q(in_s2[2]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[3]  ( .D(\outreg_stage2/N6 ), .CK(clk2), .Q(in_s2[3]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[4]  ( .D(\outreg_stage2/N7 ), .CK(clk2), .Q(in_s2[4]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[5]  ( .D(\outreg_stage2/N8 ), .CK(clk2), .Q(in_s2[5]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[6]  ( .D(\outreg_stage2/N9 ), .CK(clk2), .Q(in_s2[6]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[7]  ( .D(\outreg_stage2/N10 ), .CK(
        clk2), .Q(in_s2[7]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[8]  ( .D(\outreg_stage2/N11 ), .CK(
        clk2), .Q(in_s2[8]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[9]  ( .D(\outreg_stage2/N12 ), .CK(
        clk2), .Q(in_s2[9]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[10]  ( .D(\outreg_stage2/N13 ), .CK(
        clk2), .Q(in_s2[10]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[11]  ( .D(\outreg_stage2/N14 ), .CK(
        clk2), .Q(in_s2[11]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[12]  ( .D(\outreg_stage2/N15 ), .CK(
        clk2), .Q(in_s2[12]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[13]  ( .D(\outreg_stage2/N16 ), .CK(
        clk2), .Q(in_s2[13]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[15]  ( .D(\outreg_stage2/N18 ), .CK(
        clk2), .Q(in_s2[15]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[16]  ( .D(\outreg_stage2/N19 ), .CK(
        clk2), .Q(in_s2[16]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[17]  ( .D(\outreg_stage2/N20 ), .CK(
        clk2), .Q(in_s2[17]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[18]  ( .D(\outreg_stage2/N21 ), .CK(
        clk2), .Q(in_s2[18]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[19]  ( .D(\outreg_stage2/N22 ), .CK(
        clk2), .Q(in_s2[19]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[20]  ( .D(\outreg_stage2/N23 ), .CK(
        clk2), .Q(in_s2[20]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[21]  ( .D(\outreg_stage2/N24 ), .CK(
        clk2), .Q(in_s2[21]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[22]  ( .D(\outreg_stage2/N25 ), .CK(
        clk2), .Q(in_s2[22]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[23]  ( .D(\outreg_stage2/N26 ), .CK(
        clk2), .Q(in_s2[23]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[24]  ( .D(\outreg_stage2/N27 ), .CK(
        clk2), .Q(in_s2[24]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[25]  ( .D(\outreg_stage2/N28 ), .CK(
        clk2), .Q(in_s2[25]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[26]  ( .D(\outreg_stage2/N29 ), .CK(
        clk2), .Q(in_s2[26]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[27]  ( .D(\outreg_stage2/N30 ), .CK(
        clk2), .Q(in_s2[27]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[28]  ( .D(\outreg_stage2/N31 ), .CK(
        clk2), .Q(in_s2[28]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[30]  ( .D(\outreg_stage2/N33 ), .CK(
        clk2), .Q(in_s2[30]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[0]  ( .D(\accreg_stage2/N3 ), .CK(clk2), .Q(acc_s2[0]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[0]  ( .D(\outreg_stage2/N3 ), .CK(clk2), .Q(in_s2[0]) );
  DFFQ_X0P5M_A12TR \outreg_stage2/q_reg[31]  ( .D(\outreg_stage2/N34 ), .CK(
        clk2), .Q(in_s2[31]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[24]  ( .D(\areg_stage1/N27 ), .CK(clk1), 
        .Q(a_s1[24]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[27]  ( .D(\areg_stage1/N30 ), .CK(clk1), 
        .Q(a_s1[27]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[4]  ( .D(\areg_stage1/N7 ), .CK(clk1), 
        .Q(a_s1[4]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[7]  ( .D(\areg_stage1/N10 ), .CK(clk1), 
        .Q(a_s1[7]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[10]  ( .D(\areg_stage1/N13 ), .CK(clk1), 
        .Q(a_s1[10]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[13]  ( .D(\areg_stage1/N16 ), .CK(clk1), 
        .Q(a_s1[13]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[15]  ( .D(\areg_stage1/N18 ), .CK(clk1), 
        .Q(a_s1[15]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[21]  ( .D(\areg_stage1/N24 ), .CK(clk1), 
        .Q(a_s1[21]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[18]  ( .D(\areg_stage1/N21 ), .CK(clk1), 
        .Q(a_s1[18]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[31]  ( .D(\breg_stage1/N34 ), .CK(clk1), 
        .Q(b_s1[31]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[30]  ( .D(\areg_stage1/N33 ), .CK(clk1), 
        .Q(a_s1[30]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[1]  ( .D(\accreg_stage2/N4 ), .CK(clk2), .Q(acc_s2[1]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[2]  ( .D(\accreg_stage2/N5 ), .CK(clk2), .Q(acc_s2[2]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[3]  ( .D(\accreg_stage2/N6 ), .CK(clk2), .Q(acc_s2[3]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[4]  ( .D(\accreg_stage2/N7 ), .CK(clk2), .Q(acc_s2[4]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[5]  ( .D(\accreg_stage2/N8 ), .CK(clk2), .Q(acc_s2[5]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[6]  ( .D(\accreg_stage2/N9 ), .CK(clk2), .Q(acc_s2[6]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[7]  ( .D(\accreg_stage2/N10 ), .CK(
        clk2), .Q(acc_s2[7]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[8]  ( .D(\accreg_stage2/N11 ), .CK(
        clk2), .Q(acc_s2[8]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[9]  ( .D(\accreg_stage2/N12 ), .CK(
        clk2), .Q(acc_s2[9]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[10]  ( .D(\accreg_stage2/N13 ), .CK(
        clk2), .Q(acc_s2[10]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[11]  ( .D(\accreg_stage2/N14 ), .CK(
        clk2), .Q(acc_s2[11]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[12]  ( .D(\accreg_stage2/N15 ), .CK(
        clk2), .Q(acc_s2[12]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[13]  ( .D(\accreg_stage2/N16 ), .CK(
        clk2), .Q(acc_s2[13]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[15]  ( .D(\accreg_stage2/N18 ), .CK(
        clk2), .Q(acc_s2[15]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[16]  ( .D(\accreg_stage2/N19 ), .CK(
        clk2), .Q(acc_s2[16]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[17]  ( .D(\accreg_stage2/N20 ), .CK(
        clk2), .Q(acc_s2[17]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[18]  ( .D(\accreg_stage2/N21 ), .CK(
        clk2), .Q(acc_s2[18]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[19]  ( .D(\accreg_stage2/N22 ), .CK(
        clk2), .Q(acc_s2[19]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[20]  ( .D(\accreg_stage2/N23 ), .CK(
        clk2), .Q(acc_s2[20]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[21]  ( .D(\accreg_stage2/N24 ), .CK(
        clk2), .Q(acc_s2[21]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[22]  ( .D(\accreg_stage2/N25 ), .CK(
        clk2), .Q(acc_s2[22]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[23]  ( .D(\accreg_stage2/N26 ), .CK(
        clk2), .Q(acc_s2[23]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[24]  ( .D(\accreg_stage2/N27 ), .CK(
        clk2), .Q(acc_s2[24]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[25]  ( .D(\accreg_stage2/N28 ), .CK(
        clk2), .Q(acc_s2[25]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[26]  ( .D(\accreg_stage2/N29 ), .CK(
        clk2), .Q(acc_s2[26]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[27]  ( .D(\accreg_stage2/N30 ), .CK(
        clk2), .Q(acc_s2[27]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[28]  ( .D(\accreg_stage2/N31 ), .CK(
        clk2), .Q(acc_s2[28]) );
  DFFQ_X0P5M_A12TR \accreg_stage2/q_reg[30]  ( .D(\accreg_stage2/N33 ), .CK(
        clk2), .Q(acc_s2[30]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[12]  ( .D(\areg_stage1/N15 ), .CK(clk1), 
        .Q(a_s1[12]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[16]  ( .D(\areg_stage1/N19 ), .CK(clk1), 
        .Q(a_s1[16]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[25]  ( .D(\areg_stage1/N28 ), .CK(clk1), 
        .Q(a_s1[25]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[28]  ( .D(\areg_stage1/N31 ), .CK(clk1), 
        .Q(a_s1[28]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[9]  ( .D(\areg_stage1/N12 ), .CK(clk1), 
        .Q(a_s1[9]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[3]  ( .D(\areg_stage1/N6 ), .CK(clk1), 
        .Q(a_s1[3]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[6]  ( .D(\areg_stage1/N9 ), .CK(clk1), 
        .Q(a_s1[6]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[22]  ( .D(\areg_stage1/N25 ), .CK(clk1), 
        .Q(a_s1[22]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[19]  ( .D(\areg_stage1/N22 ), .CK(clk1), 
        .Q(a_s1[19]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[0]  ( .D(\areg_stage1/N3 ), .CK(clk1), 
        .Q(a_s1[0]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[1]  ( .D(\areg_stage1/N4 ), .CK(clk1), 
        .Q(a_s1[1]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[23]  ( .D(\areg_stage1/N26 ), .CK(clk1), 
        .Q(a_s1[23]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[30]  ( .D(\breg_stage1/N33 ), .CK(clk1), 
        .Q(b_s1[30]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[26]  ( .D(\areg_stage1/N29 ), .CK(clk1), 
        .Q(a_s1[26]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[20]  ( .D(\areg_stage1/N23 ), .CK(clk1), 
        .Q(a_s1[20]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[29]  ( .D(\breg_stage1/N32 ), .CK(clk1), 
        .Q(b_s1[29]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[28]  ( .D(\breg_stage1/N31 ), .CK(clk1), 
        .Q(b_s1[28]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[27]  ( .D(\breg_stage1/N30 ), .CK(clk1), 
        .Q(b_s1[27]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[26]  ( .D(\breg_stage1/N29 ), .CK(clk1), 
        .Q(b_s1[26]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[25]  ( .D(\breg_stage1/N28 ), .CK(clk1), 
        .Q(b_s1[25]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[23]  ( .D(\breg_stage1/N26 ), .CK(clk1), 
        .Q(b_s1[23]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[24]  ( .D(\breg_stage1/N27 ), .CK(clk1), 
        .Q(b_s1[24]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[22]  ( .D(\breg_stage1/N25 ), .CK(clk1), 
        .Q(b_s1[22]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[20]  ( .D(\breg_stage1/N23 ), .CK(clk1), 
        .Q(b_s1[20]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[21]  ( .D(\breg_stage1/N24 ), .CK(clk1), 
        .Q(b_s1[21]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[19]  ( .D(\breg_stage1/N22 ), .CK(clk1), 
        .Q(b_s1[19]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[18]  ( .D(\breg_stage1/N21 ), .CK(clk1), 
        .Q(b_s1[18]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[16]  ( .D(\breg_stage1/N19 ), .CK(clk1), 
        .Q(b_s1[16]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[17]  ( .D(\areg_stage1/N20 ), .CK(clk1), 
        .Q(a_s1[17]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[14]  ( .D(\breg_stage1/N17 ), .CK(clk1), 
        .Q(b_s1[14]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[15]  ( .D(\breg_stage1/N18 ), .CK(clk1), 
        .Q(b_s1[15]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[13]  ( .D(\breg_stage1/N16 ), .CK(clk1), 
        .Q(b_s1[13]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[12]  ( .D(\breg_stage1/N15 ), .CK(clk1), 
        .Q(b_s1[12]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[14]  ( .D(\areg_stage1/N17 ), .CK(clk1), 
        .Q(a_s1[14]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[11]  ( .D(\breg_stage1/N14 ), .CK(clk1), 
        .Q(b_s1[11]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[10]  ( .D(\breg_stage1/N13 ), .CK(clk1), 
        .Q(b_s1[10]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[8]  ( .D(\areg_stage1/N11 ), .CK(clk1), 
        .Q(a_s1[8]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[11]  ( .D(\areg_stage1/N14 ), .CK(clk1), 
        .Q(a_s1[11]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[9]  ( .D(\breg_stage1/N12 ), .CK(clk1), 
        .Q(b_s1[9]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[8]  ( .D(\breg_stage1/N11 ), .CK(clk1), 
        .Q(b_s1[8]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[7]  ( .D(\breg_stage1/N10 ), .CK(clk1), 
        .Q(b_s1[7]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[6]  ( .D(\breg_stage1/N9 ), .CK(clk1), 
        .Q(b_s1[6]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[4]  ( .D(\breg_stage1/N7 ), .CK(clk1), 
        .Q(b_s1[4]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[5]  ( .D(\breg_stage1/N8 ), .CK(clk1), 
        .Q(b_s1[5]) );
  DFFQ_X0P5M_A12TR \areg_stage1/q_reg[5]  ( .D(\areg_stage1/N8 ), .CK(clk1), 
        .Q(a_s1[5]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[2]  ( .D(\breg_stage1/N5 ), .CK(clk1), 
        .Q(b_s1[2]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[0]  ( .D(\breg_stage1/N3 ), .CK(clk1), 
        .Q(b_s1[0]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[3]  ( .D(\breg_stage1/N6 ), .CK(clk1), 
        .Q(b_s1[3]) );
  DFFQ_X0P5M_A12TR \breg_stage1/q_reg[1]  ( .D(\breg_stage1/N4 ), .CK(clk1), 
        .Q(b_s1[1]) );
  NOR2XB_X0P5M_A12TR U130 ( .BN(out[31]), .A(reset), .Y(\accreg_stage2/N34 )
         );
  NOR2XB_X0P5M_A12TR U131 ( .BN(out[30]), .A(reset), .Y(\accreg_stage2/N33 )
         );
  XOR3_X0P5M_A12TR U132 ( .A(n1272), .B(in_s2[31]), .C(acc_s2[31]), .Y(out[31]) );
  NOR2XB_X0P5M_A12TR U133 ( .BN(out[29]), .A(reset), .Y(\accreg_stage2/N32 )
         );
  NOR2XB_X0P5M_A12TR U134 ( .BN(out[28]), .A(reset), .Y(\accreg_stage2/N31 )
         );
  NOR2XB_X0P5M_A12TR U135 ( .BN(out[27]), .A(reset), .Y(\accreg_stage2/N30 )
         );
  NOR2XB_X0P5M_A12TR U136 ( .BN(out[26]), .A(reset), .Y(\accreg_stage2/N29 )
         );
  NOR2XB_X0P5M_A12TR U137 ( .BN(out[25]), .A(reset), .Y(\accreg_stage2/N28 )
         );
  NOR2XB_X0P5M_A12TR U138 ( .BN(out[24]), .A(reset), .Y(\accreg_stage2/N27 )
         );
  NOR2XB_X0P5M_A12TR U139 ( .BN(out[23]), .A(reset), .Y(\accreg_stage2/N26 )
         );
  NOR2XB_X0P5M_A12TR U140 ( .BN(out[22]), .A(reset), .Y(\accreg_stage2/N25 )
         );
  OAI222_X0P5M_A12TR U141 ( .A0(n1078), .A1(n1324), .B0(n1078), .B1(b_s1[18]), 
        .C0(n1205), .C1(n1221), .Y(n1079) );
  NOR2XB_X0P5M_A12TR U142 ( .BN(out[21]), .A(reset), .Y(\accreg_stage2/N24 )
         );
  NOR2XB_X0P5M_A12TR U143 ( .BN(out[20]), .A(reset), .Y(\accreg_stage2/N23 )
         );
  OAI222_X0P5M_A12TR U144 ( .A0(n1009), .A1(n1324), .B0(n1009), .B1(b_s1[17]), 
        .C0(n1205), .C1(n1217), .Y(n1010) );
  NOR2XB_X0P5M_A12TR U145 ( .BN(out[19]), .A(reset), .Y(\accreg_stage2/N22 )
         );
  OAI222_X0P5M_A12TR U146 ( .A0(n956), .A1(n1324), .B0(n956), .B1(b_s1[16]), 
        .C0(n1205), .C1(n1086), .Y(n957) );
  OAI222_X0P5M_A12TR U147 ( .A0(n876), .A1(n1324), .B0(n876), .B1(b_s1[15]), 
        .C0(n1205), .C1(n1237), .Y(n877) );
  NOR2XB_X0P5M_A12TR U148 ( .BN(out[18]), .A(reset), .Y(\accreg_stage2/N21 )
         );
  OAI222_X0P5M_A12TR U149 ( .A0(n814), .A1(n1324), .B0(n814), .B1(b_s1[14]), 
        .C0(n1205), .C1(n1235), .Y(n815) );
  NOR2XB_X0P5M_A12TR U150 ( .BN(out[17]), .A(reset), .Y(\accreg_stage2/N20 )
         );
  OAI222_X0P5M_A12TR U151 ( .A0(n1239), .A1(n1337), .B0(n1239), .B1(b_s1[15]), 
        .C0(n1238), .C1(n1237), .Y(n1240) );
  NOR2XB_X0P5M_A12TR U152 ( .BN(out[16]), .A(reset), .Y(\accreg_stage2/N19 )
         );
  OAI222_X0P5M_A12TR U153 ( .A0(n767), .A1(n1324), .B0(n767), .B1(b_s1[13]), 
        .C0(n1205), .C1(n1098), .Y(n768) );
  OAI222_X0P5M_A12TR U154 ( .A0(n694), .A1(n1324), .B0(n694), .B1(b_s1[12]), 
        .C0(n1205), .C1(n1025), .Y(n695) );
  OAI222_X0P5M_A12TR U155 ( .A0(n1099), .A1(n1337), .B0(n1099), .B1(b_s1[14]), 
        .C0(n1238), .C1(n1235), .Y(n1100) );
  NOR2XB_X0P5M_A12TR U156 ( .BN(out[15]), .A(reset), .Y(\accreg_stage2/N18 )
         );
  OAI222_X0P5M_A12TR U157 ( .A0(n640), .A1(n1324), .B0(n640), .B1(b_s1[11]), 
        .C0(n1205), .C1(n971), .Y(n641) );
  OAI222_X0P5M_A12TR U158 ( .A0(n1026), .A1(n1337), .B0(n1026), .B1(b_s1[13]), 
        .C0(n1238), .C1(n1098), .Y(n1027) );
  NOR2XB_X0P5M_A12TR U159 ( .BN(out[14]), .A(reset), .Y(\accreg_stage2/N17 )
         );
  OAI222_X0P5M_A12TR U160 ( .A0(n972), .A1(n1337), .B0(n972), .B1(b_s1[12]), 
        .C0(n1238), .C1(n1025), .Y(n973) );
  NOR2XB_X0P5M_A12TR U161 ( .BN(out[13]), .A(reset), .Y(\accreg_stage2/N16 )
         );
  OAI222_X0P5M_A12TR U162 ( .A0(n599), .A1(n1324), .B0(n599), .B1(b_s1[10]), 
        .C0(n1205), .C1(n892), .Y(n600) );
  NOR2XB_X0P5M_A12TR U163 ( .BN(out[12]), .A(reset), .Y(\accreg_stage2/N15 )
         );
  OAI222_X0P5M_A12TR U164 ( .A0(n893), .A1(n1337), .B0(n893), .B1(b_s1[11]), 
        .C0(n1238), .C1(n971), .Y(n894) );
  OAI222_X0P5M_A12TR U165 ( .A0(n531), .A1(n1324), .B0(n531), .B1(b_s1[9]), 
        .C0(n1205), .C1(n829), .Y(n532) );
  OAI222_X0P5M_A12TR U166 ( .A0(n482), .A1(n1324), .B0(n482), .B1(b_s1[8]), 
        .C0(n1205), .C1(n782), .Y(n483) );
  AOI211_X0P5M_A12TR U167 ( .A0(n1292), .A1(n1291), .B0(reset), .C0(n1290), 
        .Y(\outreg_stage2/N8 ) );
  NOR2XB_X0P5M_A12TR U168 ( .BN(out[11]), .A(reset), .Y(\accreg_stage2/N14 )
         );
  OAI222_X0P5M_A12TR U169 ( .A0(n830), .A1(n1337), .B0(n830), .B1(b_s1[10]), 
        .C0(n1238), .C1(n892), .Y(n831) );
  OAI222_X0P5M_A12TR U170 ( .A0(n783), .A1(n1337), .B0(n783), .B1(b_s1[9]), 
        .C0(n1238), .C1(n829), .Y(n784) );
  OAI222_X0P5M_A12TR U171 ( .A0(n445), .A1(n1324), .B0(n445), .B1(b_s1[7]), 
        .C0(n1205), .C1(n709), .Y(n446) );
  OAI222_X0P5M_A12TR U172 ( .A0(n606), .A1(n1307), .B0(n606), .B1(b_s1[9]), 
        .C0(n1222), .C1(n829), .Y(n607) );
  NOR2XB_X0P5M_A12TR U173 ( .BN(out[10]), .A(reset), .Y(\accreg_stage2/N13 )
         );
  AOI211_X0P5M_A12TR U174 ( .A0(n1287), .A1(n1286), .B0(reset), .C0(n1285), 
        .Y(\outreg_stage2/N7 ) );
  AOI211_X0P5M_A12TR U175 ( .A0(n1282), .A1(n1281), .B0(reset), .C0(n1280), 
        .Y(\outreg_stage2/N6 ) );
  OAI222_X0P5M_A12TR U176 ( .A0(n710), .A1(n1337), .B0(n710), .B1(b_s1[8]), 
        .C0(n1238), .C1(n782), .Y(n711) );
  OAI222_X0P5M_A12TR U177 ( .A0(n382), .A1(n1324), .B0(n382), .B1(b_s1[6]), 
        .C0(n1205), .C1(n655), .Y(n383) );
  OAI222_X0P5M_A12TR U178 ( .A0(n538), .A1(n1307), .B0(n538), .B1(b_s1[8]), 
        .C0(n1222), .C1(n782), .Y(n539) );
  NOR2XB_X0P5M_A12TR U179 ( .BN(out[9]), .A(reset), .Y(\accreg_stage2/N12 ) );
  OAI222_X0P5M_A12TR U180 ( .A0(n342), .A1(n1324), .B0(n342), .B1(b_s1[5]), 
        .C0(n1205), .C1(n614), .Y(n343) );
  OAI222_X0P5M_A12TR U181 ( .A0(n656), .A1(n1337), .B0(n656), .B1(b_s1[7]), 
        .C0(n1238), .C1(n709), .Y(n657) );
  NOR2XB_X0P5M_A12TR U182 ( .BN(out[8]), .A(reset), .Y(\accreg_stage2/N11 ) );
  OAI222_X0P5M_A12TR U183 ( .A0(n489), .A1(n1307), .B0(n489), .B1(b_s1[7]), 
        .C0(n1222), .C1(n709), .Y(n490) );
  OAI222_X0P5M_A12TR U184 ( .A0(n316), .A1(n1324), .B0(n316), .B1(b_s1[4]), 
        .C0(n1205), .C1(n546), .Y(n317) );
  OAI222_X0P5M_A12TR U185 ( .A0(n615), .A1(n1337), .B0(n615), .B1(b_s1[6]), 
        .C0(n1238), .C1(n655), .Y(n616) );
  OAI222_X0P5M_A12TR U186 ( .A0(n452), .A1(n1307), .B0(n452), .B1(b_s1[6]), 
        .C0(n1222), .C1(n655), .Y(n453) );
  OAI222_X0P5M_A12TR U187 ( .A0(n114), .A1(n1299), .B0(n114), .B1(b_s1[4]), 
        .C0(n1173), .C1(n546), .Y(n115) );
  NOR2XB_X0P5M_A12TR U188 ( .BN(out[7]), .A(reset), .Y(\accreg_stage2/N10 ) );
  OAI222_X0P5M_A12TR U189 ( .A0(n204), .A1(n1358), .B0(n204), .B1(b_s1[4]), 
        .C0(n1189), .C1(n546), .Y(n205) );
  OAI222_X0P5M_A12TR U190 ( .A0(n161), .A1(n1358), .B0(n161), .B1(b_s1[3]), 
        .C0(n1189), .C1(n496), .Y(n162) );
  OAI222_X0P5M_A12TR U191 ( .A0(n264), .A1(n1324), .B0(n264), .B1(b_s1[3]), 
        .C0(n1205), .C1(n496), .Y(n265) );
  NOR2XB_X0P5M_A12TR U192 ( .BN(out[6]), .A(reset), .Y(\accreg_stage2/N9 ) );
  OAI222_X0P5M_A12TR U193 ( .A0(n76), .A1(n1299), .B0(n76), .B1(b_s1[3]), .C0(
        n1173), .C1(n496), .Y(n77) );
  OAI222_X0P5M_A12TR U194 ( .A0(n389), .A1(n1307), .B0(n389), .B1(b_s1[5]), 
        .C0(n1222), .C1(n614), .Y(n390) );
  OAI222_X0P5M_A12TR U195 ( .A0(n547), .A1(n1337), .B0(n547), .B1(b_s1[5]), 
        .C0(n1238), .C1(n614), .Y(n548) );
  OAI222_X0P5M_A12TR U196 ( .A0(n134), .A1(n1358), .B0(n134), .B1(b_s1[2]), 
        .C0(n1189), .C1(n458), .Y(n135) );
  OAI222_X0P5M_A12TR U197 ( .A0(n58), .A1(n1299), .B0(n58), .B1(b_s1[2]), .C0(
        n1173), .C1(n458), .Y(n59) );
  NOR2XB_X0P5M_A12TR U198 ( .BN(out[5]), .A(reset), .Y(\accreg_stage2/N8 ) );
  OAI222_X0P5M_A12TR U199 ( .A0(n231), .A1(n1324), .B0(n231), .B1(b_s1[2]), 
        .C0(n1205), .C1(n458), .Y(n232) );
  OAI222_X0P5M_A12TR U200 ( .A0(n497), .A1(n1337), .B0(n497), .B1(b_s1[4]), 
        .C0(n1238), .C1(n546), .Y(n498) );
  OAI222_X0P5M_A12TR U201 ( .A0(n399), .A1(n1336), .B0(n399), .B1(b_s1[0]), 
        .C0(n455), .C1(n1247), .Y(n400) );
  OAI222_X0P5M_A12TR U202 ( .A0(n348), .A1(n1307), .B0(n348), .B1(b_s1[4]), 
        .C0(n1222), .C1(n546), .Y(n349) );
  OAI222_X0P5M_A12TR U203 ( .A0(n272), .A1(n1307), .B0(n272), .B1(b_s1[2]), 
        .C0(n1222), .C1(n458), .Y(n273) );
  OAI222_X0P5M_A12TR U204 ( .A0(n45), .A1(n1301), .B0(n45), .B1(n1243), .C0(
        n56), .C1(n456), .Y(n46) );
  OAI222_X0P5M_A12TR U205 ( .A0(n33), .A1(n1301), .B0(n33), .B1(n1109), .C0(
        n56), .C1(n392), .Y(n34) );
  NOR2XB_X0P5M_A12TR U206 ( .BN(out[4]), .A(reset), .Y(\accreg_stage2/N7 ) );
  OAI222_X0P5M_A12TR U207 ( .A0(n208), .A1(n1325), .B0(n208), .B1(n1243), .C0(
        n229), .C1(n456), .Y(n209) );
  OAI222_X0P5M_A12TR U208 ( .A0(n167), .A1(n1325), .B0(n167), .B1(n1109), .C0(
        n229), .C1(n392), .Y(n168) );
  OAI222_X0P5M_A12TR U209 ( .A0(n460), .A1(n1337), .B0(n460), .B1(b_s1[3]), 
        .C0(n1238), .C1(n496), .Y(n461) );
  OAI222_X0P5M_A12TR U210 ( .A0(n118), .A1(n1359), .B0(n118), .B1(n1243), .C0(
        n132), .C1(n456), .Y(n119) );
  OAI222_X0P5M_A12TR U211 ( .A0(n83), .A1(n1359), .B0(n83), .B1(n1109), .C0(
        n132), .C1(n392), .Y(n84) );
  OAI222_X0P5M_A12TR U212 ( .A0(n320), .A1(n1307), .B0(n320), .B1(b_s1[3]), 
        .C0(n1222), .C1(n496), .Y(n321) );
  AOI222_X0P5M_A12TR U213 ( .A0(a_s1[31]), .A1(n1295), .B0(a_s1[31]), .B1(
        a_s1[30]), .C0(n1295), .C1(n1294), .Y(n1296) );
  NOR2XB_X0P5M_A12TR U214 ( .BN(out[3]), .A(reset), .Y(\accreg_stage2/N6 ) );
  NOR2XB_X0P5M_A12TR U215 ( .BN(out[2]), .A(reset), .Y(\accreg_stage2/N5 ) );
  NOR2XB_X0P5M_A12TR U216 ( .BN(out[0]), .A(reset), .Y(\accreg_stage2/N3 ) );
  NOR2XB_X0P5M_A12TR U217 ( .BN(out[1]), .A(reset), .Y(\accreg_stage2/N4 ) );
  OAI22BB_X0P5M_A12TR U218 ( .A0(n1423), .A1(a_s1[6]), .B0N(a_s1[6]), .B1N(
        n1423), .Y(n79) );
  OAI22BB_X0P5M_A12TR U219 ( .A0(n1424), .A1(a_s1[22]), .B0N(a_s1[22]), .B1N(
        n1424), .Y(n717) );
  OA1B2_X0P7M_A12TR U220 ( .B0(acc_s2[0]), .B1(in_s2[0]), .A0N(n1455), .Y(
        out[0]) );
  AOI22BB_X0P5M_A12TR U221 ( .A0(a_s1[27]), .A1(n1420), .B0N(n1420), .B1N(
        a_s1[27]), .Y(n1107) );
  OAI22BB_X0P5M_A12TR U222 ( .A0(n1425), .A1(a_s1[3]), .B0N(a_s1[3]), .B1N(
        n1425), .Y(n29) );
  OAI22BB_X0P5M_A12TR U223 ( .A0(n1419), .A1(a_s1[30]), .B0N(a_s1[30]), .B1N(
        n1419), .Y(n1297) );
  AOI22BB_X0P5M_A12TR U224 ( .A0(a_s1[9]), .A1(n1384), .B0N(n1384), .B1N(
        a_s1[9]), .Y(n171) );
  OAI22BB_X0P5M_A12TR U225 ( .A0(a_s1[19]), .A1(a_s1[20]), .B0N(a_s1[20]), 
        .B1N(a_s1[19]), .Y(n550) );
  AOI22BB_X0P5M_A12TR U226 ( .A0(a_s1[17]), .A1(a_s1[18]), .B0N(a_s1[18]), 
        .B1N(a_s1[17]), .Y(n551) );
  OAI22BB_X0P5M_A12TR U227 ( .A0(a_s1[25]), .A1(a_s1[26]), .B0N(a_s1[26]), 
        .B1N(a_s1[25]), .Y(n833) );
  AOI22BB_X0P5M_A12TR U228 ( .A0(a_s1[14]), .A1(a_s1[15]), .B0N(a_s1[15]), 
        .B1N(a_s1[14]), .Y(n351) );
  OAI22BB_X0P5M_A12TR U229 ( .A0(a_s1[16]), .A1(a_s1[17]), .B0N(a_s1[17]), 
        .B1N(a_s1[16]), .Y(n396) );
  AOI22BB_X0P5M_A12TR U230 ( .A0(a_s1[8]), .A1(a_s1[7]), .B0N(a_s1[7]), .B1N(
        a_s1[8]), .Y(n81) );
  AOI22BB_X0P5M_A12TR U231 ( .A0(a_s1[11]), .A1(a_s1[10]), .B0N(a_s1[10]), 
        .B1N(a_s1[11]), .Y(n164) );
  AND2_X0P5M_A12TR U232 ( .A(acc_s2[0]), .B(in_s2[0]), .Y(n1455) );
  OAI22BB_X0P5M_A12TR U233 ( .A0(a_s1[28]), .A1(a_s1[29]), .B0N(a_s1[29]), 
        .B1N(a_s1[28]), .Y(n1106) );
  OAI22BB_X0P5M_A12TR U234 ( .A0(a_s1[12]), .A1(a_s1[11]), .B0N(a_s1[11]), 
        .B1N(a_s1[12]), .Y(n269) );
  AOI22BB_X0P5M_A12TR U235 ( .A0(a_s1[5]), .A1(a_s1[4]), .B0N(a_s1[4]), .B1N(
        a_s1[5]), .Y(n31) );
  AOI22BB_X0P5M_A12TR U236 ( .A0(a_s1[20]), .A1(a_s1[21]), .B0N(a_s1[21]), 
        .B1N(a_s1[20]), .Y(n715) );
  AOI22BB_X0P5M_A12TR U237 ( .A0(a_s1[24]), .A1(a_s1[23]), .B0N(a_s1[23]), 
        .B1N(a_s1[24]), .Y(n898) );
  AOI22BB_X0P5M_A12TR U238 ( .A0(a_s1[14]), .A1(a_s1[13]), .B0N(a_s1[13]), 
        .B1N(a_s1[14]), .Y(n267) );
  NOR2XB_X0P5M_A12TR U239 ( .BN(b[3]), .A(reset), .Y(\breg_stage1/N6 ) );
  NOR2XB_X0P5M_A12TR U240 ( .BN(a[31]), .A(reset), .Y(\areg_stage1/N34 ) );
  NOR2XB_X0P5M_A12TR U241 ( .BN(b[31]), .A(reset), .Y(\breg_stage1/N34 ) );
  NOR2XB_X0P5M_A12TR U242 ( .BN(a[18]), .A(reset), .Y(\areg_stage1/N21 ) );
  NOR2XB_X0P5M_A12TR U243 ( .BN(a[21]), .A(reset), .Y(\areg_stage1/N24 ) );
  NOR2XB_X0P5M_A12TR U244 ( .BN(a[15]), .A(reset), .Y(\areg_stage1/N18 ) );
  NOR2XB_X0P5M_A12TR U245 ( .BN(a[13]), .A(reset), .Y(\areg_stage1/N16 ) );
  NOR2XB_X0P5M_A12TR U246 ( .BN(b[1]), .A(reset), .Y(\breg_stage1/N4 ) );
  NOR2XB_X0P5M_A12TR U247 ( .BN(a[10]), .A(reset), .Y(\areg_stage1/N13 ) );
  NOR2XB_X0P5M_A12TR U248 ( .BN(a[7]), .A(reset), .Y(\areg_stage1/N10 ) );
  NOR2XB_X0P5M_A12TR U249 ( .BN(a[4]), .A(reset), .Y(\areg_stage1/N7 ) );
  NOR2XB_X0P5M_A12TR U250 ( .BN(a[27]), .A(reset), .Y(\areg_stage1/N30 ) );
  NOR2XB_X0P5M_A12TR U251 ( .BN(a[24]), .A(reset), .Y(\areg_stage1/N27 ) );
  NOR2XB_X0P5M_A12TR U252 ( .BN(a[12]), .A(reset), .Y(\areg_stage1/N15 ) );
  NOR2XB_X0P5M_A12TR U253 ( .BN(a[16]), .A(reset), .Y(\areg_stage1/N19 ) );
  NOR2XB_X0P5M_A12TR U254 ( .BN(a[25]), .A(reset), .Y(\areg_stage1/N28 ) );
  NOR2XB_X0P5M_A12TR U255 ( .BN(a[28]), .A(reset), .Y(\areg_stage1/N31 ) );
  NOR2XB_X0P5M_A12TR U256 ( .BN(a[9]), .A(reset), .Y(\areg_stage1/N12 ) );
  NOR2XB_X0P5M_A12TR U257 ( .BN(a[3]), .A(reset), .Y(\areg_stage1/N6 ) );
  NOR2XB_X0P5M_A12TR U258 ( .BN(a[6]), .A(reset), .Y(\areg_stage1/N9 ) );
  NOR2XB_X0P5M_A12TR U259 ( .BN(a[22]), .A(reset), .Y(\areg_stage1/N25 ) );
  NOR2XB_X0P5M_A12TR U260 ( .BN(a[19]), .A(reset), .Y(\areg_stage1/N22 ) );
  NOR2XB_X0P5M_A12TR U261 ( .BN(a[0]), .A(reset), .Y(\areg_stage1/N3 ) );
  NOR2XB_X0P5M_A12TR U262 ( .BN(a[1]), .A(reset), .Y(\areg_stage1/N4 ) );
  NOR2XB_X0P5M_A12TR U263 ( .BN(a[23]), .A(reset), .Y(\areg_stage1/N26 ) );
  NOR2XB_X0P5M_A12TR U264 ( .BN(b[30]), .A(reset), .Y(\breg_stage1/N33 ) );
  NOR2XB_X0P5M_A12TR U265 ( .BN(a[26]), .A(reset), .Y(\areg_stage1/N29 ) );
  NOR2XB_X0P5M_A12TR U266 ( .BN(a[20]), .A(reset), .Y(\areg_stage1/N23 ) );
  NOR2XB_X0P5M_A12TR U267 ( .BN(b[29]), .A(reset), .Y(\breg_stage1/N32 ) );
  NOR2XB_X0P5M_A12TR U268 ( .BN(b[28]), .A(reset), .Y(\breg_stage1/N31 ) );
  NOR2XB_X0P5M_A12TR U269 ( .BN(b[27]), .A(reset), .Y(\breg_stage1/N30 ) );
  NOR2XB_X0P5M_A12TR U270 ( .BN(b[26]), .A(reset), .Y(\breg_stage1/N29 ) );
  NOR2XB_X0P5M_A12TR U271 ( .BN(b[25]), .A(reset), .Y(\breg_stage1/N28 ) );
  NOR2XB_X0P5M_A12TR U272 ( .BN(b[23]), .A(reset), .Y(\breg_stage1/N26 ) );
  NOR2XB_X0P5M_A12TR U273 ( .BN(b[24]), .A(reset), .Y(\breg_stage1/N27 ) );
  NOR2XB_X0P5M_A12TR U274 ( .BN(b[22]), .A(reset), .Y(\breg_stage1/N25 ) );
  NOR2XB_X0P5M_A12TR U275 ( .BN(b[20]), .A(reset), .Y(\breg_stage1/N23 ) );
  NOR2XB_X0P5M_A12TR U276 ( .BN(b[21]), .A(reset), .Y(\breg_stage1/N24 ) );
  NOR2XB_X0P5M_A12TR U277 ( .BN(b[19]), .A(reset), .Y(\breg_stage1/N22 ) );
  NOR2XB_X0P5M_A12TR U278 ( .BN(b[18]), .A(reset), .Y(\breg_stage1/N21 ) );
  NOR2XB_X0P5M_A12TR U279 ( .BN(b[17]), .A(reset), .Y(\breg_stage1/N20 ) );
  NOR2XB_X0P5M_A12TR U280 ( .BN(a[30]), .A(reset), .Y(\areg_stage1/N33 ) );
  NOR2XB_X0P5M_A12TR U281 ( .BN(b[12]), .A(reset), .Y(\breg_stage1/N15 ) );
  NOR2XB_X0P5M_A12TR U282 ( .BN(b[6]), .A(reset), .Y(\breg_stage1/N9 ) );
  NOR2XB_X0P5M_A12TR U283 ( .BN(a[29]), .A(reset), .Y(\areg_stage1/N32 ) );
  NOR2XB_X0P5M_A12TR U284 ( .BN(b[7]), .A(reset), .Y(\breg_stage1/N10 ) );
  NOR2XB_X0P5M_A12TR U285 ( .BN(b[16]), .A(reset), .Y(\breg_stage1/N19 ) );
  NOR2XB_X0P5M_A12TR U286 ( .BN(a[2]), .A(reset), .Y(\areg_stage1/N5 ) );
  NOR2XB_X0P5M_A12TR U287 ( .BN(b[15]), .A(reset), .Y(\breg_stage1/N18 ) );
  NOR2XB_X0P5M_A12TR U288 ( .BN(a[5]), .A(reset), .Y(\areg_stage1/N8 ) );
  NOR2XB_X0P5M_A12TR U289 ( .BN(a[17]), .A(reset), .Y(\areg_stage1/N20 ) );
  NOR2XB_X0P5M_A12TR U290 ( .BN(b[11]), .A(reset), .Y(\breg_stage1/N14 ) );
  NOR2XB_X0P5M_A12TR U291 ( .BN(b[14]), .A(reset), .Y(\breg_stage1/N17 ) );
  NOR2XB_X0P5M_A12TR U292 ( .BN(b[2]), .A(reset), .Y(\breg_stage1/N5 ) );
  NOR2XB_X0P5M_A12TR U293 ( .BN(b[10]), .A(reset), .Y(\breg_stage1/N13 ) );
  NOR2XB_X0P5M_A12TR U294 ( .BN(b[0]), .A(reset), .Y(\breg_stage1/N3 ) );
  NOR2XB_X0P5M_A12TR U295 ( .BN(a[8]), .A(reset), .Y(\areg_stage1/N11 ) );
  NOR2XB_X0P5M_A12TR U296 ( .BN(b[9]), .A(reset), .Y(\breg_stage1/N12 ) );
  NOR2XB_X0P5M_A12TR U297 ( .BN(a[14]), .A(reset), .Y(\areg_stage1/N17 ) );
  NOR2XB_X0P5M_A12TR U298 ( .BN(a[11]), .A(reset), .Y(\areg_stage1/N14 ) );
  NOR2XB_X0P5M_A12TR U299 ( .BN(b[4]), .A(reset), .Y(\breg_stage1/N7 ) );
  NOR2XB_X0P5M_A12TR U300 ( .BN(b[8]), .A(reset), .Y(\breg_stage1/N11 ) );
  NOR2XB_X0P5M_A12TR U301 ( .BN(b[13]), .A(reset), .Y(\breg_stage1/N16 ) );
  NOR2XB_X0P5M_A12TR U302 ( .BN(b[5]), .A(reset), .Y(\breg_stage1/N8 ) );
  INV_X0P5B_A12TR U303 ( .A(a_s1[2]), .Y(n1425) );
  INV_X0P5B_A12TR U304 ( .A(a_s1[0]), .Y(n2) );
  NAND2_X0P5A_A12TR U305 ( .A(n2), .B(a_s1[1]), .Y(n1370) );
  INV_X0P5B_A12TR U306 ( .A(n1370), .Y(n22) );
  NAND2_X0P5A_A12TR U307 ( .A(n1425), .B(n22), .Y(n28) );
  INV_X0P5B_A12TR U308 ( .A(n28), .Y(n1162) );
  INV_X0P5B_A12TR U309 ( .A(b_s1[2]), .Y(n458) );
  INV_X0P5B_A12TR U310 ( .A(b_s1[0]), .Y(n1247) );
  INV_X0P5B_A12TR U311 ( .A(b_s1[1]), .Y(n393) );
  AOI21_X0P5M_A12TR U312 ( .A0(n458), .A1(n1247), .B0(n393), .Y(n16) );
  NAND3_X0P5M_A12TR U313 ( .A(a_s1[1]), .B(a_s1[0]), .C(n1425), .Y(n15) );
  OAI31_X0P5M_A12TR U314 ( .A0(a_s1[1]), .A1(n1425), .A2(n2), .B0(n15), .Y(
        n1141) );
  INV_X0P5B_A12TR U315 ( .A(n1141), .Y(n1371) );
  INV_X0P5B_A12TR U316 ( .A(n1371), .Y(n1373) );
  INV_X0P5B_A12TR U317 ( .A(b_s1[4]), .Y(n546) );
  NOR3_X0P7M_A12TR U318 ( .A(a_s1[1]), .B(a_s1[0]), .C(n1425), .Y(n1376) );
  NOR3_X0P7M_A12TR U319 ( .A(n2), .B(a_s1[2]), .C(a_s1[1]), .Y(n1156) );
  AOI31_X0P5M_A12TR U320 ( .A0(a_s1[1]), .A1(a_s1[2]), .A2(a_s1[0]), .B0(n1156), .Y(n25) );
  INV_X0P5B_A12TR U321 ( .A(n25), .Y(n1375) );
  AOI22_X0P5M_A12TR U322 ( .A0(n1376), .A1(b_s1[3]), .B0(b_s1[5]), .B1(n1375), 
        .Y(n3) );
  OAI211_X0P5M_A12TR U323 ( .A0(n546), .A1(n1370), .B0(a_s1[2]), .C0(n3), .Y(
        n5) );
  INV_X0P5B_A12TR U324 ( .A(n15), .Y(n1157) );
  AOI22_X0P5M_A12TR U325 ( .A0(n1157), .A1(n1118), .B0(n1156), .B1(b_s1[5]), 
        .Y(n4) );
  AO21A1AI2_X0P5M_A12TR U326 ( .A0(n1118), .A1(n1373), .B0(n5), .C0(n4), .Y(n6) );
  AOI21_X0P5M_A12TR U327 ( .A0(n1162), .A1(b_s1[4]), .B0(n6), .Y(n1289) );
  NAND2_X0P5A_A12TR U328 ( .A(b_s1[0]), .B(n29), .Y(n38) );
  INV_X0P5B_A12TR U329 ( .A(n38), .Y(n1282) );
  INV_X0P5B_A12TR U330 ( .A(n29), .Y(n7) );
  NOR2_X0P5B_A12TR U331 ( .A(n31), .B(n7), .Y(n1302) );
  XNOR2_X0P5M_A12TR U332 ( .A(a_s1[3]), .B(a_s1[4]), .Y(n30) );
  NOR2_X0P5B_A12TR U333 ( .A(n29), .B(n30), .Y(n1303) );
  AOI22_X0P5M_A12TR U334 ( .A0(b_s1[1]), .A1(b_s1[0]), .B0(n1247), .B1(n393), 
        .Y(n1298) );
  AND2_X0P5M_A12TR U335 ( .A(n31), .B(n29), .Y(n1301) );
  AOI222_X0P5M_A12TR U336 ( .A0(b_s1[1]), .A1(n1302), .B0(b_s1[0]), .B1(n1303), 
        .C0(n1298), .C1(n1301), .Y(n36) );
  NAND3_X0P5M_A12TR U337 ( .A(a_s1[5]), .B(n1282), .C(n36), .Y(n8) );
  AO21A1AI2_X0P5M_A12TR U338 ( .A0(n1282), .A1(a_s1[5]), .B0(n36), .C0(n8), 
        .Y(n1284) );
  AOI222_X0P5M_A12TR U339 ( .A0(n1375), .A1(b_s1[1]), .B0(n22), .B1(b_s1[0]), 
        .C0(n1373), .C1(n1298), .Y(n1274) );
  NAND2_X0P5A_A12TR U340 ( .A(a_s1[2]), .B(n1274), .Y(n9) );
  AOI21_X0P5M_A12TR U341 ( .A0(a_s1[0]), .A1(b_s1[0]), .B0(n9), .Y(n1277) );
  NAND3_X0P5M_A12TR U342 ( .A(b_s1[1]), .B(n1247), .C(b_s1[2]), .Y(n10) );
  AO21A1AI2_X0P5M_A12TR U343 ( .A0(n1247), .A1(b_s1[1]), .B0(b_s1[2]), .C0(n10), .Y(n392) );
  AOI22_X0P5M_A12TR U344 ( .A0(b_s1[1]), .A1(n1162), .B0(n1156), .B1(b_s1[2]), 
        .Y(n14) );
  AOI21_X0P5M_A12TR U345 ( .A0(b_s1[1]), .A1(n22), .B0(n1425), .Y(n12) );
  AOI22_X0P5M_A12TR U346 ( .A0(n1376), .A1(b_s1[0]), .B0(b_s1[2]), .B1(n1375), 
        .Y(n11) );
  OAI211_X0P5M_A12TR U347 ( .A0(n1371), .A1(n392), .B0(n12), .C0(n11), .Y(n13)
         );
  OAI211_X0P5M_A12TR U348 ( .A0(n392), .A1(n15), .B0(n14), .C0(n13), .Y(n1276)
         );
  NAND2_X0P5A_A12TR U349 ( .A(n1277), .B(n1276), .Y(n1278) );
  ADDF_X1M_A12TR U350 ( .A(b_s1[2]), .B(b_s1[3]), .CI(n16), .CO(n21), .S(n1243) );
  AOI22_X0P5M_A12TR U351 ( .A0(b_s1[1]), .A1(n1376), .B0(b_s1[3]), .B1(n1375), 
        .Y(n17) );
  OAI211_X0P5M_A12TR U352 ( .A0(n1370), .A1(n458), .B0(a_s1[2]), .C0(n17), .Y(
        n19) );
  AOI22_X0P5M_A12TR U353 ( .A0(n1243), .A1(n1157), .B0(b_s1[3]), .B1(n1156), 
        .Y(n18) );
  AO21A1AI2_X0P5M_A12TR U354 ( .A0(n1243), .A1(n1373), .B0(n19), .C0(n18), .Y(
        n20) );
  AOI21_X0P5M_A12TR U355 ( .A0(b_s1[2]), .A1(n1162), .B0(n20), .Y(n1279) );
  AOI21_X0P5M_A12TR U356 ( .A0(n1278), .A1(n38), .B0(n1279), .Y(n1287) );
  INV_X0P5B_A12TR U357 ( .A(b_s1[3]), .Y(n496) );
  ADDF_X1M_A12TR U358 ( .A(b_s1[3]), .B(b_s1[4]), .CI(n21), .CO(n39), .S(n1342) );
  AOI22_X0P5M_A12TR U359 ( .A0(n1157), .A1(n1342), .B0(n1156), .B1(b_s1[4]), 
        .Y(n27) );
  AOI21_X0P5M_A12TR U360 ( .A0(b_s1[3]), .A1(n22), .B0(n1425), .Y(n24) );
  AOI22_X0P5M_A12TR U361 ( .A0(b_s1[2]), .A1(n1376), .B0(n1342), .B1(n1373), 
        .Y(n23) );
  OAI211_X0P5M_A12TR U362 ( .A0(n25), .A1(n546), .B0(n24), .C0(n23), .Y(n26)
         );
  OAI211_X0P5M_A12TR U363 ( .A0(n28), .A1(n496), .B0(n27), .C0(n26), .Y(n1283)
         );
  CGENI_X1M_A12TR U364 ( .A(n1284), .B(n1287), .CI(n1283), .CON(n1292) );
  INV_X0P5B_A12TR U365 ( .A(a_s1[5]), .Y(n1423) );
  NOR3BB_X0P5M_A12TR U366 ( .AN(n31), .BN(n30), .C(n29), .Y(n1299) );
  NAND2_X0P5A_A12TR U367 ( .A(n1423), .B(n1299), .Y(n1173) );
  INV_X0P5B_A12TR U368 ( .A(n1173), .Y(n48) );
  NAND2_X0P5A_A12TR U369 ( .A(n1303), .B(n1423), .Y(n1168) );
  NAND2_X0P5A_A12TR U370 ( .A(n1302), .B(n1423), .Y(n1167) );
  OAI22_X0P5M_A12TR U371 ( .A0(n393), .A1(n1168), .B0(n458), .B1(n1167), .Y(
        n35) );
  INV_X0P5B_A12TR U372 ( .A(n1303), .Y(n1170) );
  AOI22_X0P5M_A12TR U373 ( .A0(b_s1[2]), .A1(n1302), .B0(b_s1[0]), .B1(n1299), 
        .Y(n32) );
  OAI211_X0P5M_A12TR U374 ( .A0(n393), .A1(n1170), .B0(a_s1[5]), .C0(n32), .Y(
        n33) );
  INV_X0P5B_A12TR U375 ( .A(n392), .Y(n1109) );
  NAND2_X0P5A_A12TR U376 ( .A(n1301), .B(n1423), .Y(n56) );
  AOI211_X0P5M_A12TR U377 ( .A0(b_s1[0]), .A1(n48), .B0(n35), .C0(n34), .Y(n54) );
  AND2_X0P5M_A12TR U378 ( .A(n36), .B(a_s1[5]), .Y(n37) );
  NAND2_X0P5A_A12TR U379 ( .A(n38), .B(n37), .Y(n53) );
  XNOR2_X0P5M_A12TR U380 ( .A(n54), .B(n53), .Y(n1288) );
  CGEN_X1M_A12TR U381 ( .A(n1289), .B(n1292), .CI(n1288), .CO(n69) );
  ADDF_X1M_A12TR U382 ( .A(b_s1[4]), .B(b_s1[5]), .CI(n39), .CO(n62), .S(n1118) );
  INV_X0P5B_A12TR U383 ( .A(b_s1[5]), .Y(n614) );
  AOI22_X0P5M_A12TR U384 ( .A0(n1376), .A1(b_s1[4]), .B0(b_s1[6]), .B1(n1375), 
        .Y(n40) );
  OAI211_X0P5M_A12TR U385 ( .A0(n614), .A1(n1370), .B0(a_s1[2]), .C0(n40), .Y(
        n42) );
  AOI22_X0P5M_A12TR U386 ( .A0(n1157), .A1(n1253), .B0(n1156), .B1(b_s1[6]), 
        .Y(n41) );
  AO21A1AI2_X0P5M_A12TR U387 ( .A0(n1253), .A1(n1373), .B0(n42), .C0(n41), .Y(
        n43) );
  AOI21_X0P5M_A12TR U388 ( .A0(n1162), .A1(b_s1[5]), .B0(n43), .Y(n68) );
  NAND2_X0P5A_A12TR U389 ( .A(b_s1[0]), .B(n79), .Y(n88) );
  OAI22_X0P5M_A12TR U390 ( .A0(n496), .A1(n1167), .B0(n458), .B1(n1168), .Y(
        n47) );
  AOI22_X0P5M_A12TR U391 ( .A0(b_s1[1]), .A1(n1299), .B0(b_s1[3]), .B1(n1302), 
        .Y(n44) );
  OAI211_X0P5M_A12TR U392 ( .A0(n458), .A1(n1170), .B0(a_s1[5]), .C0(n44), .Y(
        n45) );
  INV_X0P5B_A12TR U393 ( .A(n1243), .Y(n456) );
  AOI211_X0P5M_A12TR U394 ( .A0(b_s1[1]), .A1(n48), .B0(n47), .C0(n46), .Y(n52) );
  OAI21_X0P5M_A12TR U395 ( .A0(n54), .A1(n53), .B0(n52), .Y(n49) );
  OAI31_X0P5M_A12TR U396 ( .A0(n54), .A1(n52), .A2(n53), .B0(n49), .Y(n50) );
  XNOR2_X0P5M_A12TR U397 ( .A(n88), .B(n50), .Y(n67) );
  NOR2_X0P5B_A12TR U398 ( .A(reset), .B(n51), .Y(\outreg_stage2/N9 ) );
  OA21A1OI2_X0P7M_A12TR U399 ( .A0(n54), .A1(n53), .B0(n88), .C0(n52), .Y(n55)
         );
  INV_X0P5B_A12TR U400 ( .A(n55), .Y(n74) );
  INV_X0P5B_A12TR U401 ( .A(n56), .Y(n1178) );
  OAI22_X0P5M_A12TR U402 ( .A0(n496), .A1(n1168), .B0(n546), .B1(n1167), .Y(
        n60) );
  AOI22_X0P5M_A12TR U403 ( .A0(n1301), .A1(n1342), .B0(n1302), .B1(b_s1[4]), 
        .Y(n57) );
  OAI211_X0P5M_A12TR U404 ( .A0(n496), .A1(n1170), .B0(a_s1[5]), .C0(n57), .Y(
        n58) );
  AOI211_X0P5M_A12TR U405 ( .A0(n1342), .A1(n1178), .B0(n60), .C0(n59), .Y(n73) );
  INV_X0P5B_A12TR U406 ( .A(a_s1[8]), .Y(n1384) );
  NOR2_X0P5B_A12TR U407 ( .A(n1384), .B(n88), .Y(n61) );
  AND2_X0P5M_A12TR U408 ( .A(n79), .B(n81), .Y(n1359) );
  NOR2XB_X0P5M_A12TR U409 ( .BN(n79), .A(n81), .Y(n1362) );
  XNOR2_X0P5M_A12TR U410 ( .A(a_s1[6]), .B(a_s1[7]), .Y(n80) );
  NOR2_X0P5B_A12TR U411 ( .A(n79), .B(n80), .Y(n1361) );
  AOI222_X0P5M_A12TR U412 ( .A0(n1359), .A1(n1298), .B0(n1362), .B1(b_s1[1]), 
        .C0(b_s1[0]), .C1(n1361), .Y(n86) );
  XOR2_X0P5M_A12TR U413 ( .A(n61), .B(n86), .Y(n72) );
  ADDF_X1M_A12TR U414 ( .A(b_s1[5]), .B(b_s1[6]), .CI(n62), .CO(n91), .S(n1253) );
  INV_X0P5B_A12TR U415 ( .A(b_s1[6]), .Y(n655) );
  AOI22_X0P5M_A12TR U416 ( .A0(n1376), .A1(b_s1[5]), .B0(b_s1[7]), .B1(n1375), 
        .Y(n63) );
  OAI211_X0P5M_A12TR U417 ( .A0(n655), .A1(n1370), .B0(a_s1[2]), .C0(n63), .Y(
        n65) );
  AOI22_X0P5M_A12TR U418 ( .A0(n1157), .A1(n1378), .B0(n1156), .B1(b_s1[7]), 
        .Y(n64) );
  AO21A1AI2_X0P5M_A12TR U419 ( .A0(n1378), .A1(n1373), .B0(n65), .C0(n64), .Y(
        n66) );
  AOI21_X0P5M_A12TR U420 ( .A0(n1162), .A1(b_s1[6]), .B0(n66), .Y(n97) );
  ADDF_X1M_A12TR U421 ( .A(n69), .B(n68), .CI(n67), .CO(n96), .S(n51) );
  XNOR2_X0P5M_A12TR U422 ( .A(n97), .B(n96), .Y(n71) );
  INV_X0P5B_A12TR U423 ( .A(reset), .Y(n1450) );
  OAI21_X0P5M_A12TR U424 ( .A0(n98), .A1(n71), .B0(n1450), .Y(n70) );
  AOI21_X0P5M_A12TR U425 ( .A0(n98), .A1(n71), .B0(n70), .Y(
        \outreg_stage2/N10 ) );
  ADDF_X1M_A12TR U426 ( .A(n74), .B(n73), .CI(n72), .CO(n112), .S(n98) );
  OAI22_X0P5M_A12TR U427 ( .A0(n546), .A1(n1168), .B0(n614), .B1(n1167), .Y(
        n78) );
  AOI22_X0P5M_A12TR U428 ( .A0(n1301), .A1(n1118), .B0(n1302), .B1(b_s1[5]), 
        .Y(n75) );
  OAI211_X0P5M_A12TR U429 ( .A0(n546), .A1(n1170), .B0(a_s1[5]), .C0(n75), .Y(
        n76) );
  AOI211_X0P5M_A12TR U430 ( .A0(n1118), .A1(n1178), .B0(n78), .C0(n77), .Y(
        n111) );
  NOR3BB_X0P5M_A12TR U431 ( .AN(n81), .BN(n80), .C(n79), .Y(n1358) );
  NAND2_X0P5A_A12TR U432 ( .A(n1384), .B(n1358), .Y(n1189) );
  INV_X0P5B_A12TR U433 ( .A(n1189), .Y(n121) );
  NAND2_X0P5A_A12TR U434 ( .A(n1361), .B(n1384), .Y(n1184) );
  NAND2_X0P5A_A12TR U435 ( .A(n1362), .B(n1384), .Y(n1182) );
  OAI22_X0P5M_A12TR U436 ( .A0(n393), .A1(n1184), .B0(n458), .B1(n1182), .Y(
        n85) );
  INV_X0P5B_A12TR U437 ( .A(n1361), .Y(n1187) );
  AOI22_X0P5M_A12TR U438 ( .A0(b_s1[2]), .A1(n1362), .B0(b_s1[0]), .B1(n1358), 
        .Y(n82) );
  OAI211_X0P5M_A12TR U439 ( .A0(n393), .A1(n1187), .B0(a_s1[8]), .C0(n82), .Y(
        n83) );
  NAND2_X0P5A_A12TR U440 ( .A(n1359), .B(n1384), .Y(n132) );
  AOI211_X0P5M_A12TR U441 ( .A0(b_s1[0]), .A1(n121), .B0(n85), .C0(n84), .Y(
        n90) );
  AND2_X0P5M_A12TR U442 ( .A(n86), .B(a_s1[8]), .Y(n87) );
  NAND2_X0P5A_A12TR U443 ( .A(n88), .B(n87), .Y(n89) );
  NOR2_X0P5B_A12TR U444 ( .A(n90), .B(n89), .Y(n131) );
  AO21_X0P5M_A12TR U445 ( .A0(n90), .A1(n89), .B0(n131), .Y(n110) );
  ADDF_X1M_A12TR U446 ( .A(b_s1[6]), .B(b_s1[7]), .CI(n91), .CO(n105), .S(
        n1378) );
  INV_X0P5B_A12TR U447 ( .A(b_s1[7]), .Y(n709) );
  AOI22_X0P5M_A12TR U448 ( .A0(n1376), .A1(b_s1[6]), .B0(b_s1[8]), .B1(n1375), 
        .Y(n92) );
  OAI211_X0P5M_A12TR U449 ( .A0(n709), .A1(n1370), .B0(a_s1[2]), .C0(n92), .Y(
        n94) );
  AOI22_X0P5M_A12TR U450 ( .A0(n1157), .A1(n1125), .B0(n1156), .B1(b_s1[8]), 
        .Y(n93) );
  AO21A1AI2_X0P5M_A12TR U451 ( .A0(n1125), .A1(n1141), .B0(n94), .C0(n93), .Y(
        n95) );
  AOI21_X0P5M_A12TR U452 ( .A0(n1162), .A1(b_s1[7]), .B0(n95), .Y(n102) );
  XOR2_X0P5M_A12TR U453 ( .A(n103), .B(n102), .Y(n100) );
  CGENI_X1M_A12TR U454 ( .A(n98), .B(n97), .CI(n96), .CON(n101) );
  OAI21_X0P5M_A12TR U455 ( .A0(n100), .A1(n101), .B0(n1450), .Y(n99) );
  AOI21_X0P5M_A12TR U456 ( .A0(n100), .A1(n101), .B0(n99), .Y(
        \outreg_stage2/N11 ) );
  INV_X0P5B_A12TR U457 ( .A(n101), .Y(n104) );
  CGEN_X1M_A12TR U458 ( .A(n104), .B(n103), .CI(n102), .CO(n147) );
  ADDF_X1M_A12TR U459 ( .A(b_s1[7]), .B(b_s1[8]), .CI(n105), .CO(n140), .S(
        n1125) );
  INV_X0P5B_A12TR U460 ( .A(b_s1[8]), .Y(n782) );
  AOI22_X0P5M_A12TR U461 ( .A0(n1376), .A1(b_s1[7]), .B0(b_s1[9]), .B1(n1375), 
        .Y(n106) );
  OAI211_X0P5M_A12TR U462 ( .A0(n782), .A1(n1370), .B0(a_s1[2]), .C0(n106), 
        .Y(n108) );
  AOI22_X0P5M_A12TR U463 ( .A0(n1157), .A1(n1260), .B0(n1156), .B1(b_s1[9]), 
        .Y(n107) );
  AO21A1AI2_X0P5M_A12TR U464 ( .A0(n1260), .A1(n1141), .B0(n108), .C0(n107), 
        .Y(n109) );
  AOI21_X0P5M_A12TR U465 ( .A0(n1162), .A1(b_s1[8]), .B0(n109), .Y(n146) );
  ADDF_X1M_A12TR U466 ( .A(n112), .B(n111), .CI(n110), .CO(n125), .S(n103) );
  OAI22_X0P5M_A12TR U467 ( .A0(n614), .A1(n1168), .B0(n1167), .B1(n655), .Y(
        n116) );
  AOI22_X0P5M_A12TR U468 ( .A0(n1301), .A1(n1253), .B0(n1302), .B1(b_s1[6]), 
        .Y(n113) );
  OAI211_X0P5M_A12TR U469 ( .A0(n614), .A1(n1170), .B0(a_s1[5]), .C0(n113), 
        .Y(n114) );
  AOI211_X0P5M_A12TR U470 ( .A0(n1178), .A1(n1253), .B0(n116), .C0(n115), .Y(
        n124) );
  OAI22_X0P5M_A12TR U471 ( .A0(n496), .A1(n1182), .B0(n458), .B1(n1184), .Y(
        n120) );
  AOI22_X0P5M_A12TR U472 ( .A0(b_s1[1]), .A1(n1358), .B0(b_s1[3]), .B1(n1362), 
        .Y(n117) );
  OAI211_X0P5M_A12TR U473 ( .A0(n458), .A1(n1187), .B0(a_s1[8]), .C0(n117), 
        .Y(n118) );
  AOI211_X0P5M_A12TR U474 ( .A0(b_s1[1]), .A1(n121), .B0(n120), .C0(n119), .Y(
        n130) );
  NOR2_X0P5B_A12TR U475 ( .A(n1247), .B(n171), .Y(n139) );
  XOR3_X0P5M_A12TR U476 ( .A(n131), .B(n130), .C(n139), .Y(n123) );
  NOR2_X0P5B_A12TR U477 ( .A(reset), .B(n122), .Y(\outreg_stage2/N12 ) );
  ADDF_X1M_A12TR U478 ( .A(n125), .B(n124), .CI(n123), .CO(n152), .S(n145) );
  OAI22_X0P5M_A12TR U479 ( .A0(n1168), .A1(n655), .B0(n1167), .B1(n709), .Y(
        n129) );
  AOI22_X0P5M_A12TR U480 ( .A0(n1301), .A1(n1378), .B0(n1302), .B1(b_s1[7]), 
        .Y(n126) );
  OAI211_X0P5M_A12TR U481 ( .A0(n655), .A1(n1170), .B0(a_s1[5]), .C0(n126), 
        .Y(n127) );
  OAI222_X0P5M_A12TR U482 ( .A0(n127), .A1(n1299), .B0(n127), .B1(b_s1[5]), 
        .C0(n1173), .C1(n614), .Y(n128) );
  AOI211_X0P5M_A12TR U483 ( .A0(n1178), .A1(n1378), .B0(n129), .C0(n128), .Y(
        n151) );
  OAI21B_X0P5M_A12TR U484 ( .A0(n139), .A1(n131), .B0N(n130), .Y(n159) );
  INV_X0P5B_A12TR U485 ( .A(n132), .Y(n1194) );
  OAI22_X0P5M_A12TR U486 ( .A0(n496), .A1(n1184), .B0(n546), .B1(n1182), .Y(
        n136) );
  AOI22_X0P5M_A12TR U487 ( .A0(n1342), .A1(n1359), .B0(b_s1[4]), .B1(n1362), 
        .Y(n133) );
  OAI211_X0P5M_A12TR U488 ( .A0(n496), .A1(n1187), .B0(a_s1[8]), .C0(n133), 
        .Y(n134) );
  AOI211_X0P5M_A12TR U489 ( .A0(n1342), .A1(n1194), .B0(n136), .C0(n135), .Y(
        n158) );
  NOR2XB_X0P5M_A12TR U490 ( .BN(n164), .A(n171), .Y(n1325) );
  NOR2_X0P5B_A12TR U491 ( .A(n164), .B(n171), .Y(n1328) );
  XNOR2_X0P5M_A12TR U492 ( .A(a_s1[9]), .B(a_s1[10]), .Y(n165) );
  NAND2XB_X0P5M_A12TR U493 ( .BN(n165), .A(n171), .Y(n1203) );
  INV_X0P5B_A12TR U494 ( .A(n1203), .Y(n1327) );
  AOI222_X0P5M_A12TR U495 ( .A0(n1325), .A1(n1298), .B0(n1328), .B1(b_s1[1]), 
        .C0(b_s1[0]), .C1(n1327), .Y(n137) );
  INV_X0P5B_A12TR U496 ( .A(n137), .Y(n170) );
  NAND3_X0P5M_A12TR U497 ( .A(n139), .B(a_s1[11]), .C(n170), .Y(n138) );
  AO21A1AI2_X0P5M_A12TR U498 ( .A0(a_s1[11]), .A1(n139), .B0(n170), .C0(n138), 
        .Y(n157) );
  ADDF_X1M_A12TR U499 ( .A(b_s1[8]), .B(b_s1[9]), .CI(n140), .CO(n174), .S(
        n1260) );
  INV_X0P5B_A12TR U500 ( .A(b_s1[9]), .Y(n829) );
  AOI22_X0P5M_A12TR U501 ( .A0(n1376), .A1(b_s1[8]), .B0(b_s1[10]), .B1(n1375), 
        .Y(n141) );
  OAI211_X0P5M_A12TR U502 ( .A0(n829), .A1(n1370), .B0(a_s1[2]), .C0(n141), 
        .Y(n143) );
  AOI22_X0P5M_A12TR U503 ( .A0(n1157), .A1(n1332), .B0(n1156), .B1(b_s1[10]), 
        .Y(n142) );
  AO21A1AI2_X0P5M_A12TR U504 ( .A0(n1332), .A1(n1141), .B0(n143), .C0(n142), 
        .Y(n144) );
  AOI21_X0P5M_A12TR U505 ( .A0(n1162), .A1(b_s1[9]), .B0(n144), .Y(n180) );
  ADDF_X1M_A12TR U506 ( .A(n147), .B(n146), .CI(n145), .CO(n179), .S(n122) );
  XNOR2_X0P5M_A12TR U507 ( .A(n180), .B(n179), .Y(n149) );
  OAI21_X0P5M_A12TR U508 ( .A0(n181), .A1(n149), .B0(n1450), .Y(n148) );
  AOI21_X0P5M_A12TR U509 ( .A0(n181), .A1(n149), .B0(n148), .Y(
        \outreg_stage2/N13 ) );
  ADDF_X1M_A12TR U510 ( .A(n152), .B(n151), .CI(n150), .CO(n195), .S(n181) );
  OAI22_X0P5M_A12TR U511 ( .A0(n1168), .A1(n709), .B0(n1167), .B1(n782), .Y(
        n156) );
  AOI22_X0P5M_A12TR U512 ( .A0(n1301), .A1(n1125), .B0(n1302), .B1(b_s1[8]), 
        .Y(n153) );
  OAI211_X0P5M_A12TR U513 ( .A0(n709), .A1(n1170), .B0(a_s1[5]), .C0(n153), 
        .Y(n154) );
  OAI222_X0P5M_A12TR U514 ( .A0(n154), .A1(n1299), .B0(n154), .B1(b_s1[6]), 
        .C0(n1173), .C1(n655), .Y(n155) );
  AOI211_X0P5M_A12TR U515 ( .A0(n1178), .A1(n1125), .B0(n156), .C0(n155), .Y(
        n194) );
  ADDF_X1M_A12TR U516 ( .A(n159), .B(n158), .CI(n157), .CO(n202), .S(n150) );
  OAI22_X0P5M_A12TR U517 ( .A0(n546), .A1(n1184), .B0(n614), .B1(n1182), .Y(
        n163) );
  AOI22_X0P5M_A12TR U518 ( .A0(n1118), .A1(n1359), .B0(b_s1[5]), .B1(n1362), 
        .Y(n160) );
  OAI211_X0P5M_A12TR U519 ( .A0(n546), .A1(n1187), .B0(a_s1[8]), .C0(n160), 
        .Y(n161) );
  AOI211_X0P5M_A12TR U520 ( .A0(n1118), .A1(n1194), .B0(n163), .C0(n162), .Y(
        n201) );
  INV_X0P5B_A12TR U521 ( .A(a_s1[11]), .Y(n1426) );
  AND3_X0P5M_A12TR U522 ( .A(n171), .B(n165), .C(n164), .Y(n1324) );
  NAND2_X0P5A_A12TR U523 ( .A(n1426), .B(n1324), .Y(n1205) );
  INV_X0P5B_A12TR U524 ( .A(n1205), .Y(n211) );
  NAND2_X0P5A_A12TR U525 ( .A(n1327), .B(n1426), .Y(n1200) );
  NAND2_X0P5A_A12TR U526 ( .A(n1328), .B(n1426), .Y(n1198) );
  OAI22_X0P5M_A12TR U527 ( .A0(n393), .A1(n1200), .B0(n458), .B1(n1198), .Y(
        n169) );
  AOI22_X0P5M_A12TR U528 ( .A0(b_s1[2]), .A1(n1328), .B0(b_s1[0]), .B1(n1324), 
        .Y(n166) );
  OAI211_X0P5M_A12TR U529 ( .A0(n393), .A1(n1203), .B0(a_s1[11]), .C0(n166), 
        .Y(n167) );
  NAND2_X0P5A_A12TR U530 ( .A(n1325), .B(n1426), .Y(n229) );
  AOI211_X0P5M_A12TR U531 ( .A0(b_s1[0]), .A1(n211), .B0(n169), .C0(n168), .Y(
        n173) );
  OAI211_X0P5M_A12TR U532 ( .A0(n1247), .A1(n171), .B0(a_s1[11]), .C0(n137), 
        .Y(n172) );
  NOR2_X0P5B_A12TR U533 ( .A(n173), .B(n172), .Y(n228) );
  AO21_X0P5M_A12TR U534 ( .A0(n173), .A1(n172), .B0(n228), .Y(n200) );
  ADDF_X1M_A12TR U535 ( .A(b_s1[9]), .B(b_s1[10]), .CI(n174), .CO(n188), .S(
        n1332) );
  INV_X0P5B_A12TR U536 ( .A(b_s1[10]), .Y(n892) );
  AOI22_X0P5M_A12TR U537 ( .A0(n1376), .A1(b_s1[9]), .B0(b_s1[11]), .B1(n1375), 
        .Y(n175) );
  OAI211_X0P5M_A12TR U538 ( .A0(n892), .A1(n1370), .B0(a_s1[2]), .C0(n175), 
        .Y(n177) );
  AOI22_X0P5M_A12TR U539 ( .A0(n1157), .A1(n1132), .B0(n1156), .B1(b_s1[11]), 
        .Y(n176) );
  AO21A1AI2_X0P5M_A12TR U540 ( .A0(n1132), .A1(n1141), .B0(n177), .C0(n176), 
        .Y(n178) );
  AOI21_X0P5M_A12TR U541 ( .A0(n1162), .A1(b_s1[10]), .B0(n178), .Y(n185) );
  XOR2_X0P5M_A12TR U542 ( .A(n186), .B(n185), .Y(n183) );
  CGENI_X1M_A12TR U543 ( .A(n181), .B(n180), .CI(n179), .CON(n184) );
  OAI21_X0P5M_A12TR U544 ( .A0(n183), .A1(n184), .B0(n1450), .Y(n182) );
  AOI21_X0P5M_A12TR U545 ( .A0(n183), .A1(n184), .B0(n182), .Y(
        \outreg_stage2/N14 ) );
  INV_X0P5B_A12TR U546 ( .A(n184), .Y(n187) );
  CGEN_X1M_A12TR U547 ( .A(n187), .B(n186), .CI(n185), .CO(n243) );
  ADDF_X1M_A12TR U548 ( .A(b_s1[10]), .B(b_s1[11]), .CI(n188), .CO(n236), .S(
        n1132) );
  INV_X0P5B_A12TR U549 ( .A(b_s1[11]), .Y(n971) );
  AOI22_X0P5M_A12TR U550 ( .A0(n1376), .A1(b_s1[10]), .B0(b_s1[12]), .B1(n1375), .Y(n189) );
  OAI211_X0P5M_A12TR U551 ( .A0(n971), .A1(n1370), .B0(a_s1[2]), .C0(n189), 
        .Y(n191) );
  AOI22_X0P5M_A12TR U552 ( .A0(n1157), .A1(n1267), .B0(n1156), .B1(b_s1[12]), 
        .Y(n190) );
  AO21A1AI2_X0P5M_A12TR U553 ( .A0(n1267), .A1(n1141), .B0(n191), .C0(n190), 
        .Y(n192) );
  AOI21_X0P5M_A12TR U554 ( .A0(n1162), .A1(b_s1[11]), .B0(n192), .Y(n242) );
  ADDF_X1M_A12TR U555 ( .A(n195), .B(n194), .CI(n193), .CO(n215), .S(n186) );
  OAI22_X0P5M_A12TR U556 ( .A0(n1168), .A1(n782), .B0(n1167), .B1(n829), .Y(
        n199) );
  AOI22_X0P5M_A12TR U557 ( .A0(n1301), .A1(n1260), .B0(n1302), .B1(b_s1[9]), 
        .Y(n196) );
  OAI211_X0P5M_A12TR U558 ( .A0(n782), .A1(n1170), .B0(a_s1[5]), .C0(n196), 
        .Y(n197) );
  OAI222_X0P5M_A12TR U559 ( .A0(n197), .A1(n1299), .B0(n197), .B1(b_s1[7]), 
        .C0(n1173), .C1(n709), .Y(n198) );
  AOI211_X0P5M_A12TR U560 ( .A0(n1178), .A1(n1260), .B0(n199), .C0(n198), .Y(
        n214) );
  ADDF_X1M_A12TR U561 ( .A(n202), .B(n201), .CI(n200), .CO(n222), .S(n193) );
  OAI22_X0P5M_A12TR U562 ( .A0(n614), .A1(n1184), .B0(n655), .B1(n1182), .Y(
        n206) );
  AOI22_X0P5M_A12TR U563 ( .A0(b_s1[6]), .A1(n1362), .B0(n1359), .B1(n1253), 
        .Y(n203) );
  OAI211_X0P5M_A12TR U564 ( .A0(n614), .A1(n1187), .B0(a_s1[8]), .C0(n203), 
        .Y(n204) );
  AOI211_X0P5M_A12TR U565 ( .A0(n1194), .A1(n1253), .B0(n206), .C0(n205), .Y(
        n221) );
  OAI22_X0P5M_A12TR U566 ( .A0(n496), .A1(n1198), .B0(n458), .B1(n1200), .Y(
        n210) );
  AOI22_X0P5M_A12TR U567 ( .A0(b_s1[1]), .A1(n1324), .B0(b_s1[3]), .B1(n1328), 
        .Y(n207) );
  OAI211_X0P5M_A12TR U568 ( .A0(n458), .A1(n1203), .B0(a_s1[11]), .C0(n207), 
        .Y(n208) );
  AOI211_X0P5M_A12TR U569 ( .A0(b_s1[1]), .A1(n211), .B0(n210), .C0(n209), .Y(
        n227) );
  NOR2_X0P5B_A12TR U570 ( .A(n1247), .B(n269), .Y(n276) );
  XOR3_X0P5M_A12TR U571 ( .A(n227), .B(n228), .C(n276), .Y(n220) );
  NOR2_X0P5B_A12TR U572 ( .A(reset), .B(n212), .Y(\outreg_stage2/N15 ) );
  ADDF_X1M_A12TR U573 ( .A(n215), .B(n214), .CI(n213), .CO(n248), .S(n241) );
  OAI22_X0P5M_A12TR U574 ( .A0(n1168), .A1(n829), .B0(n1167), .B1(n892), .Y(
        n219) );
  AOI22_X0P5M_A12TR U575 ( .A0(n1301), .A1(n1332), .B0(n1302), .B1(b_s1[10]), 
        .Y(n216) );
  OAI211_X0P5M_A12TR U576 ( .A0(n829), .A1(n1170), .B0(a_s1[5]), .C0(n216), 
        .Y(n217) );
  OAI222_X0P5M_A12TR U577 ( .A0(n217), .A1(n1299), .B0(n217), .B1(b_s1[8]), 
        .C0(n1173), .C1(n782), .Y(n218) );
  AOI211_X0P5M_A12TR U578 ( .A0(n1178), .A1(n1332), .B0(n219), .C0(n218), .Y(
        n247) );
  ADDF_X1M_A12TR U579 ( .A(n222), .B(n221), .CI(n220), .CO(n255), .S(n213) );
  OAI22_X0P5M_A12TR U580 ( .A0(n655), .A1(n1184), .B0(n709), .B1(n1182), .Y(
        n226) );
  AOI22_X0P5M_A12TR U581 ( .A0(n1378), .A1(n1359), .B0(b_s1[7]), .B1(n1362), 
        .Y(n223) );
  OAI211_X0P5M_A12TR U582 ( .A0(n655), .A1(n1187), .B0(a_s1[8]), .C0(n223), 
        .Y(n224) );
  OAI222_X0P5M_A12TR U583 ( .A0(n224), .A1(n1358), .B0(n224), .B1(b_s1[5]), 
        .C0(n1189), .C1(n614), .Y(n225) );
  AOI211_X0P5M_A12TR U584 ( .A0(n1378), .A1(n1194), .B0(n226), .C0(n225), .Y(
        n254) );
  OAI21B_X0P5M_A12TR U585 ( .A0(n276), .A1(n228), .B0N(n227), .Y(n262) );
  INV_X0P5B_A12TR U586 ( .A(n229), .Y(n1210) );
  OAI22_X0P5M_A12TR U587 ( .A0(n496), .A1(n1200), .B0(n546), .B1(n1198), .Y(
        n233) );
  AOI22_X0P5M_A12TR U588 ( .A0(n1342), .A1(n1325), .B0(b_s1[4]), .B1(n1328), 
        .Y(n230) );
  OAI211_X0P5M_A12TR U589 ( .A0(n496), .A1(n1203), .B0(a_s1[11]), .C0(n230), 
        .Y(n231) );
  AOI211_X0P5M_A12TR U590 ( .A0(n1342), .A1(n1210), .B0(n233), .C0(n232), .Y(
        n261) );
  NAND2XB_X0P5M_A12TR U591 ( .BN(n269), .A(n267), .Y(n1219) );
  INV_X0P5B_A12TR U592 ( .A(n1219), .Y(n1305) );
  NOR2_X0P5B_A12TR U593 ( .A(n267), .B(n269), .Y(n1307) );
  XNOR2_X0P5M_A12TR U594 ( .A(a_s1[12]), .B(a_s1[13]), .Y(n268) );
  NAND2XB_X0P5M_A12TR U595 ( .BN(n268), .A(n269), .Y(n883) );
  INV_X0P5B_A12TR U596 ( .A(n883), .Y(n1308) );
  AOI222_X0P5M_A12TR U597 ( .A0(n1305), .A1(n1298), .B0(n1307), .B1(b_s1[1]), 
        .C0(n1308), .C1(b_s1[0]), .Y(n234) );
  INV_X0P5B_A12TR U598 ( .A(n234), .Y(n275) );
  NAND3_X0P5M_A12TR U599 ( .A(n276), .B(a_s1[14]), .C(n275), .Y(n235) );
  AO21A1AI2_X0P5M_A12TR U600 ( .A0(a_s1[14]), .A1(n276), .B0(n275), .C0(n235), 
        .Y(n260) );
  ADDF_X1M_A12TR U601 ( .A(b_s1[11]), .B(b_s1[12]), .CI(n236), .CO(n279), .S(
        n1267) );
  INV_X0P5B_A12TR U602 ( .A(b_s1[12]), .Y(n1025) );
  AOI22_X0P5M_A12TR U603 ( .A0(n1376), .A1(b_s1[11]), .B0(b_s1[13]), .B1(n1375), .Y(n237) );
  OAI211_X0P5M_A12TR U604 ( .A0(n1025), .A1(n1370), .B0(a_s1[2]), .C0(n237), 
        .Y(n239) );
  AOI22_X0P5M_A12TR U605 ( .A0(n1157), .A1(n1312), .B0(n1156), .B1(b_s1[13]), 
        .Y(n238) );
  AO21A1AI2_X0P5M_A12TR U606 ( .A0(n1312), .A1(n1373), .B0(n239), .C0(n238), 
        .Y(n240) );
  AOI21_X0P5M_A12TR U607 ( .A0(n1162), .A1(b_s1[12]), .B0(n240), .Y(n285) );
  ADDF_X1M_A12TR U608 ( .A(n243), .B(n242), .CI(n241), .CO(n284), .S(n212) );
  XNOR2_X0P5M_A12TR U609 ( .A(n285), .B(n284), .Y(n245) );
  OAI21_X0P5M_A12TR U610 ( .A0(n286), .A1(n245), .B0(n1450), .Y(n244) );
  AOI21_X0P5M_A12TR U611 ( .A0(n286), .A1(n245), .B0(n244), .Y(
        \outreg_stage2/N16 ) );
  ADDF_X1M_A12TR U612 ( .A(n248), .B(n247), .CI(n246), .CO(n300), .S(n286) );
  OAI22_X0P5M_A12TR U613 ( .A0(n1168), .A1(n892), .B0(n1167), .B1(n971), .Y(
        n252) );
  AOI22_X0P5M_A12TR U614 ( .A0(n1301), .A1(n1132), .B0(n1302), .B1(b_s1[11]), 
        .Y(n249) );
  OAI211_X0P5M_A12TR U615 ( .A0(n892), .A1(n1170), .B0(a_s1[5]), .C0(n249), 
        .Y(n250) );
  OAI222_X0P5M_A12TR U616 ( .A0(n250), .A1(n1299), .B0(n250), .B1(b_s1[9]), 
        .C0(n1173), .C1(n829), .Y(n251) );
  AOI211_X0P5M_A12TR U617 ( .A0(n1178), .A1(n1132), .B0(n252), .C0(n251), .Y(
        n299) );
  ADDF_X1M_A12TR U618 ( .A(n255), .B(n254), .CI(n253), .CO(n307), .S(n246) );
  OAI22_X0P5M_A12TR U619 ( .A0(n709), .A1(n1184), .B0(n782), .B1(n1182), .Y(
        n259) );
  AOI22_X0P5M_A12TR U620 ( .A0(n1359), .A1(n1125), .B0(n1362), .B1(b_s1[8]), 
        .Y(n256) );
  OAI211_X0P5M_A12TR U621 ( .A0(n709), .A1(n1187), .B0(a_s1[8]), .C0(n256), 
        .Y(n257) );
  OAI222_X0P5M_A12TR U622 ( .A0(n257), .A1(n1358), .B0(n257), .B1(b_s1[6]), 
        .C0(n1189), .C1(n655), .Y(n258) );
  AOI211_X0P5M_A12TR U623 ( .A0(n1194), .A1(n1125), .B0(n259), .C0(n258), .Y(
        n306) );
  ADDF_X1M_A12TR U624 ( .A(n262), .B(n261), .CI(n260), .CO(n314), .S(n253) );
  OAI22_X0P5M_A12TR U625 ( .A0(n546), .A1(n1200), .B0(n614), .B1(n1198), .Y(
        n266) );
  AOI22_X0P5M_A12TR U626 ( .A0(n1118), .A1(n1325), .B0(b_s1[5]), .B1(n1328), 
        .Y(n263) );
  OAI211_X0P5M_A12TR U627 ( .A0(n546), .A1(n1203), .B0(a_s1[11]), .C0(n263), 
        .Y(n264) );
  AOI211_X0P5M_A12TR U628 ( .A0(n1118), .A1(n1210), .B0(n266), .C0(n265), .Y(
        n313) );
  NAND3_X0P5M_A12TR U629 ( .A(n269), .B(n268), .C(n267), .Y(n270) );
  NOR2_X0P5B_A12TR U630 ( .A(a_s1[14]), .B(n270), .Y(n1226) );
  INV_X0P5B_A12TR U631 ( .A(a_s1[14]), .Y(n1385) );
  NAND2_X0P5A_A12TR U632 ( .A(n1308), .B(n1385), .Y(n1216) );
  NAND2_X0P5A_A12TR U633 ( .A(n1305), .B(n1385), .Y(n1215) );
  OAI22_X0P5M_A12TR U634 ( .A0(n393), .A1(n1216), .B0(n392), .B1(n1215), .Y(
        n274) );
  INV_X0P5B_A12TR U635 ( .A(n270), .Y(n1304) );
  AOI22_X0P5M_A12TR U636 ( .A0(b_s1[0]), .A1(n1304), .B0(n1109), .B1(n1305), 
        .Y(n271) );
  OAI211_X0P5M_A12TR U637 ( .A0(n393), .A1(n883), .B0(a_s1[14]), .C0(n271), 
        .Y(n272) );
  NAND2_X0P5A_A12TR U638 ( .A(n1307), .B(n1385), .Y(n1222) );
  AOI211_X0P5M_A12TR U639 ( .A0(b_s1[0]), .A1(n1226), .B0(n274), .C0(n273), 
        .Y(n278) );
  NAND3BB_X0P5M_A12TR U640 ( .AN(n276), .BN(n1385), .C(n234), .Y(n277) );
  NOR2_X0P5B_A12TR U641 ( .A(n278), .B(n277), .Y(n346) );
  AO21_X0P5M_A12TR U642 ( .A0(n278), .A1(n277), .B0(n346), .Y(n312) );
  ADDF_X1M_A12TR U643 ( .A(b_s1[12]), .B(b_s1[13]), .CI(n279), .CO(n293), .S(
        n1312) );
  INV_X0P5B_A12TR U644 ( .A(b_s1[13]), .Y(n1098) );
  AOI22_X0P5M_A12TR U645 ( .A0(n1376), .A1(b_s1[12]), .B0(b_s1[14]), .B1(n1375), .Y(n280) );
  OAI211_X0P5M_A12TR U646 ( .A0(n1098), .A1(n1370), .B0(a_s1[2]), .C0(n280), 
        .Y(n282) );
  AOI22_X0P5M_A12TR U647 ( .A0(n1157), .A1(n1096), .B0(n1156), .B1(b_s1[14]), 
        .Y(n281) );
  AO21A1AI2_X0P5M_A12TR U648 ( .A0(n1096), .A1(n1141), .B0(n282), .C0(n281), 
        .Y(n283) );
  AOI21_X0P5M_A12TR U649 ( .A0(n1162), .A1(b_s1[13]), .B0(n283), .Y(n290) );
  XOR2_X0P5M_A12TR U650 ( .A(n291), .B(n290), .Y(n288) );
  CGENI_X1M_A12TR U651 ( .A(n286), .B(n285), .CI(n284), .CON(n289) );
  OAI21_X0P5M_A12TR U652 ( .A0(n288), .A1(n289), .B0(n1450), .Y(n287) );
  AOI21_X0P5M_A12TR U653 ( .A0(n288), .A1(n289), .B0(n287), .Y(
        \outreg_stage2/N17 ) );
  INV_X0P5B_A12TR U654 ( .A(n289), .Y(n292) );
  CGEN_X1M_A12TR U655 ( .A(n292), .B(n291), .CI(n290), .CO(n361) );
  ADDF_X1M_A12TR U656 ( .A(b_s1[13]), .B(b_s1[14]), .CI(n293), .CO(n354), .S(
        n1096) );
  INV_X0P5B_A12TR U657 ( .A(b_s1[14]), .Y(n1235) );
  AOI22_X0P5M_A12TR U658 ( .A0(n1376), .A1(b_s1[13]), .B0(b_s1[15]), .B1(n1375), .Y(n294) );
  OAI211_X0P5M_A12TR U659 ( .A0(n1235), .A1(n1370), .B0(a_s1[2]), .C0(n294), 
        .Y(n296) );
  AOI22_X0P5M_A12TR U660 ( .A0(n1157), .A1(n1233), .B0(n1156), .B1(b_s1[15]), 
        .Y(n295) );
  AO21A1AI2_X0P5M_A12TR U661 ( .A0(n1233), .A1(n1373), .B0(n296), .C0(n295), 
        .Y(n297) );
  AOI21_X0P5M_A12TR U662 ( .A0(n1162), .A1(b_s1[14]), .B0(n297), .Y(n360) );
  ADDF_X1M_A12TR U663 ( .A(n300), .B(n299), .CI(n298), .CO(n326), .S(n291) );
  OAI22_X0P5M_A12TR U664 ( .A0(n1168), .A1(n971), .B0(n1167), .B1(n1025), .Y(
        n304) );
  AOI22_X0P5M_A12TR U665 ( .A0(n1301), .A1(n1267), .B0(n1302), .B1(b_s1[12]), 
        .Y(n301) );
  OAI211_X0P5M_A12TR U666 ( .A0(n971), .A1(n1170), .B0(a_s1[5]), .C0(n301), 
        .Y(n302) );
  OAI222_X0P5M_A12TR U667 ( .A0(n302), .A1(n1299), .B0(n302), .B1(b_s1[10]), 
        .C0(n1173), .C1(n892), .Y(n303) );
  AOI211_X0P5M_A12TR U668 ( .A0(n1178), .A1(n1267), .B0(n304), .C0(n303), .Y(
        n325) );
  ADDF_X1M_A12TR U669 ( .A(n307), .B(n306), .CI(n305), .CO(n333), .S(n298) );
  OAI22_X0P5M_A12TR U670 ( .A0(n782), .A1(n1184), .B0(n829), .B1(n1182), .Y(
        n311) );
  AOI22_X0P5M_A12TR U671 ( .A0(n1359), .A1(n1260), .B0(n1362), .B1(b_s1[9]), 
        .Y(n308) );
  OAI211_X0P5M_A12TR U672 ( .A0(n782), .A1(n1187), .B0(a_s1[8]), .C0(n308), 
        .Y(n309) );
  OAI222_X0P5M_A12TR U673 ( .A0(n309), .A1(n1358), .B0(n309), .B1(b_s1[7]), 
        .C0(n1189), .C1(n709), .Y(n310) );
  AOI211_X0P5M_A12TR U674 ( .A0(n1194), .A1(n1260), .B0(n311), .C0(n310), .Y(
        n332) );
  ADDF_X1M_A12TR U675 ( .A(n314), .B(n313), .CI(n312), .CO(n340), .S(n305) );
  OAI22_X0P5M_A12TR U676 ( .A0(n614), .A1(n1200), .B0(n655), .B1(n1198), .Y(
        n318) );
  AOI22_X0P5M_A12TR U677 ( .A0(b_s1[6]), .A1(n1328), .B0(n1325), .B1(n1253), 
        .Y(n315) );
  OAI211_X0P5M_A12TR U678 ( .A0(n614), .A1(n1203), .B0(a_s1[11]), .C0(n315), 
        .Y(n316) );
  AOI211_X0P5M_A12TR U679 ( .A0(n1210), .A1(n1253), .B0(n318), .C0(n317), .Y(
        n339) );
  OAI22_X0P5M_A12TR U680 ( .A0(n456), .A1(n1215), .B0(n458), .B1(n1216), .Y(
        n322) );
  AOI22_X0P5M_A12TR U681 ( .A0(n1243), .A1(n1305), .B0(b_s1[1]), .B1(n1304), 
        .Y(n319) );
  OAI211_X0P5M_A12TR U682 ( .A0(n458), .A1(n883), .B0(a_s1[14]), .C0(n319), 
        .Y(n320) );
  AOI211_X0P5M_A12TR U683 ( .A0(b_s1[1]), .A1(n1226), .B0(n322), .C0(n321), 
        .Y(n345) );
  INV_X0P5B_A12TR U684 ( .A(n351), .Y(n397) );
  NOR2_X0P5B_A12TR U685 ( .A(n1247), .B(n397), .Y(n402) );
  XOR3_X0P5M_A12TR U686 ( .A(n345), .B(n346), .C(n402), .Y(n338) );
  NOR2_X0P5B_A12TR U687 ( .A(reset), .B(n323), .Y(\outreg_stage2/N18 ) );
  ADDF_X1M_A12TR U688 ( .A(n326), .B(n325), .CI(n324), .CO(n366), .S(n359) );
  OAI22_X0P5M_A12TR U689 ( .A0(n1168), .A1(n1025), .B0(n1167), .B1(n1098), .Y(
        n330) );
  AOI22_X0P5M_A12TR U690 ( .A0(n1301), .A1(n1312), .B0(n1302), .B1(b_s1[13]), 
        .Y(n327) );
  OAI211_X0P5M_A12TR U691 ( .A0(n1025), .A1(n1170), .B0(a_s1[5]), .C0(n327), 
        .Y(n328) );
  OAI222_X0P5M_A12TR U692 ( .A0(n328), .A1(n1299), .B0(n328), .B1(b_s1[11]), 
        .C0(n1173), .C1(n971), .Y(n329) );
  AOI211_X0P5M_A12TR U693 ( .A0(n1178), .A1(n1312), .B0(n330), .C0(n329), .Y(
        n365) );
  ADDF_X1M_A12TR U694 ( .A(n333), .B(n332), .CI(n331), .CO(n373), .S(n324) );
  OAI22_X0P5M_A12TR U695 ( .A0(n892), .A1(n1182), .B0(n829), .B1(n1184), .Y(
        n337) );
  AOI22_X0P5M_A12TR U696 ( .A0(n1359), .A1(n1332), .B0(n1362), .B1(b_s1[10]), 
        .Y(n334) );
  OAI211_X0P5M_A12TR U697 ( .A0(n829), .A1(n1187), .B0(a_s1[8]), .C0(n334), 
        .Y(n335) );
  OAI222_X0P5M_A12TR U698 ( .A0(n335), .A1(n1358), .B0(n335), .B1(b_s1[8]), 
        .C0(n1189), .C1(n782), .Y(n336) );
  AOI211_X0P5M_A12TR U699 ( .A0(n1332), .A1(n1194), .B0(n337), .C0(n336), .Y(
        n372) );
  ADDF_X1M_A12TR U700 ( .A(n340), .B(n339), .CI(n338), .CO(n380), .S(n331) );
  OAI22_X0P5M_A12TR U701 ( .A0(n655), .A1(n1200), .B0(n709), .B1(n1198), .Y(
        n344) );
  AOI22_X0P5M_A12TR U702 ( .A0(n1378), .A1(n1325), .B0(b_s1[7]), .B1(n1328), 
        .Y(n341) );
  OAI211_X0P5M_A12TR U703 ( .A0(n655), .A1(n1203), .B0(a_s1[11]), .C0(n341), 
        .Y(n342) );
  AOI211_X0P5M_A12TR U704 ( .A0(n1378), .A1(n1210), .B0(n344), .C0(n343), .Y(
        n379) );
  OAI21B_X0P5M_A12TR U705 ( .A0(n402), .A1(n346), .B0N(n345), .Y(n387) );
  INV_X0P5B_A12TR U706 ( .A(n1342), .Y(n494) );
  OAI22_X0P5M_A12TR U707 ( .A0(n496), .A1(n1216), .B0(n494), .B1(n1215), .Y(
        n350) );
  AOI22_X0P5M_A12TR U708 ( .A0(b_s1[2]), .A1(n1304), .B0(n1342), .B1(n1305), 
        .Y(n347) );
  OAI211_X0P5M_A12TR U709 ( .A0(n496), .A1(n883), .B0(a_s1[14]), .C0(n347), 
        .Y(n348) );
  AOI211_X0P5M_A12TR U710 ( .A0(b_s1[2]), .A1(n1226), .B0(n350), .C0(n349), 
        .Y(n386) );
  NOR2_X0P5B_A12TR U711 ( .A(n396), .B(n397), .Y(n1334) );
  NAND2_X0P5A_A12TR U712 ( .A(n396), .B(n351), .Y(n395) );
  INV_X0P5B_A12TR U713 ( .A(n395), .Y(n1337) );
  XNOR2_X0P5M_A12TR U714 ( .A(a_s1[16]), .B(a_s1[15]), .Y(n398) );
  NOR2_X0P5B_A12TR U715 ( .A(n351), .B(n398), .Y(n1338) );
  AOI222_X0P5M_A12TR U716 ( .A0(n1334), .A1(n1298), .B0(n1337), .B1(b_s1[1]), 
        .C0(n1338), .C1(b_s1[0]), .Y(n352) );
  INV_X0P5B_A12TR U717 ( .A(n352), .Y(n403) );
  NAND3_X0P5M_A12TR U718 ( .A(n402), .B(a_s1[17]), .C(n403), .Y(n353) );
  AO21A1AI2_X0P5M_A12TR U719 ( .A0(a_s1[17]), .A1(n402), .B0(n403), .C0(n353), 
        .Y(n385) );
  ADDF_X1M_A12TR U720 ( .A(b_s1[14]), .B(b_s1[15]), .CI(n354), .CO(n408), .S(
        n1233) );
  INV_X0P5B_A12TR U721 ( .A(b_s1[15]), .Y(n1237) );
  AOI22_X0P5M_A12TR U722 ( .A0(n1376), .A1(b_s1[14]), .B0(b_s1[16]), .B1(n1375), .Y(n355) );
  OAI211_X0P5M_A12TR U723 ( .A0(n1237), .A1(n1370), .B0(a_s1[2]), .C0(n355), 
        .Y(n357) );
  AOI22_X0P5M_A12TR U724 ( .A0(n1157), .A1(n1335), .B0(n1156), .B1(b_s1[16]), 
        .Y(n356) );
  AO21A1AI2_X0P5M_A12TR U725 ( .A0(n1335), .A1(n1141), .B0(n357), .C0(n356), 
        .Y(n358) );
  AOI21_X0P5M_A12TR U726 ( .A0(n1162), .A1(b_s1[15]), .B0(n358), .Y(n414) );
  ADDF_X1M_A12TR U727 ( .A(n361), .B(n360), .CI(n359), .CO(n413), .S(n323) );
  XNOR2_X0P5M_A12TR U728 ( .A(n414), .B(n413), .Y(n363) );
  OAI21_X0P5M_A12TR U729 ( .A0(n415), .A1(n363), .B0(n1450), .Y(n362) );
  AOI21_X0P5M_A12TR U730 ( .A0(n415), .A1(n363), .B0(n362), .Y(
        \outreg_stage2/N19 ) );
  ADDF_X1M_A12TR U731 ( .A(n366), .B(n365), .CI(n364), .CO(n429), .S(n415) );
  OAI22_X0P5M_A12TR U732 ( .A0(n1168), .A1(n1098), .B0(n1167), .B1(n1235), .Y(
        n370) );
  AOI22_X0P5M_A12TR U733 ( .A0(n1301), .A1(n1096), .B0(n1302), .B1(b_s1[14]), 
        .Y(n367) );
  OAI211_X0P5M_A12TR U734 ( .A0(n1098), .A1(n1170), .B0(a_s1[5]), .C0(n367), 
        .Y(n368) );
  OAI222_X0P5M_A12TR U735 ( .A0(n368), .A1(n1299), .B0(n368), .B1(b_s1[12]), 
        .C0(n1173), .C1(n1025), .Y(n369) );
  AOI211_X0P5M_A12TR U736 ( .A0(n1178), .A1(n1096), .B0(n370), .C0(n369), .Y(
        n428) );
  ADDF_X1M_A12TR U737 ( .A(n373), .B(n372), .CI(n371), .CO(n436), .S(n364) );
  OAI22_X0P5M_A12TR U738 ( .A0(n971), .A1(n1182), .B0(n892), .B1(n1184), .Y(
        n377) );
  AOI22_X0P5M_A12TR U739 ( .A0(n1359), .A1(n1132), .B0(n1362), .B1(b_s1[11]), 
        .Y(n374) );
  OAI211_X0P5M_A12TR U740 ( .A0(n892), .A1(n1187), .B0(a_s1[8]), .C0(n374), 
        .Y(n375) );
  OAI222_X0P5M_A12TR U741 ( .A0(n375), .A1(n1358), .B0(n375), .B1(b_s1[9]), 
        .C0(n1189), .C1(n829), .Y(n376) );
  AOI211_X0P5M_A12TR U742 ( .A0(n1194), .A1(n1132), .B0(n377), .C0(n376), .Y(
        n435) );
  ADDF_X1M_A12TR U743 ( .A(n380), .B(n379), .CI(n378), .CO(n443), .S(n371) );
  OAI22_X0P5M_A12TR U744 ( .A0(n709), .A1(n1200), .B0(n782), .B1(n1198), .Y(
        n384) );
  AOI22_X0P5M_A12TR U745 ( .A0(n1325), .A1(n1125), .B0(n1328), .B1(b_s1[8]), 
        .Y(n381) );
  OAI211_X0P5M_A12TR U746 ( .A0(n709), .A1(n1203), .B0(a_s1[11]), .C0(n381), 
        .Y(n382) );
  AOI211_X0P5M_A12TR U747 ( .A0(n1210), .A1(n1125), .B0(n384), .C0(n383), .Y(
        n442) );
  ADDF_X1M_A12TR U748 ( .A(n387), .B(n386), .CI(n385), .CO(n450), .S(n378) );
  INV_X0P5B_A12TR U749 ( .A(n1118), .Y(n544) );
  OAI22_X0P5M_A12TR U750 ( .A0(n546), .A1(n1216), .B0(n544), .B1(n1215), .Y(
        n391) );
  AOI22_X0P5M_A12TR U751 ( .A0(b_s1[3]), .A1(n1304), .B0(n1118), .B1(n1305), 
        .Y(n388) );
  OAI211_X0P5M_A12TR U752 ( .A0(n546), .A1(n883), .B0(a_s1[14]), .C0(n388), 
        .Y(n389) );
  AOI211_X0P5M_A12TR U753 ( .A0(b_s1[3]), .A1(n1226), .B0(n391), .C0(n390), 
        .Y(n449) );
  NOR2_X0P5B_A12TR U754 ( .A(n395), .B(a_s1[17]), .Y(n459) );
  INV_X0P5B_A12TR U755 ( .A(a_s1[17]), .Y(n1382) );
  NAND2_X0P5A_A12TR U756 ( .A(n1338), .B(n1382), .Y(n1232) );
  NAND2_X0P5A_A12TR U757 ( .A(n1334), .B(n1382), .Y(n1231) );
  OAI22_X0P5M_A12TR U758 ( .A0(n393), .A1(n1232), .B0(n392), .B1(n1231), .Y(
        n401) );
  AOI22_X0P5M_A12TR U759 ( .A0(b_s1[1]), .A1(n1338), .B0(n1109), .B1(n1334), 
        .Y(n394) );
  OAI211_X0P5M_A12TR U760 ( .A0(n458), .A1(n395), .B0(a_s1[17]), .C0(n394), 
        .Y(n399) );
  NOR3BB_X0P5M_A12TR U761 ( .AN(n398), .BN(n397), .C(n396), .Y(n1336) );
  NAND2_X0P5A_A12TR U762 ( .A(n1382), .B(n1336), .Y(n455) );
  AOI211_X0P5M_A12TR U763 ( .A0(b_s1[2]), .A1(n459), .B0(n401), .C0(n400), .Y(
        n407) );
  INV_X0P5B_A12TR U764 ( .A(n402), .Y(n405) );
  NOR2_X0P5B_A12TR U765 ( .A(n1382), .B(n403), .Y(n404) );
  NAND2_X0P5A_A12TR U766 ( .A(n405), .B(n404), .Y(n406) );
  NOR2_X0P5B_A12TR U767 ( .A(n407), .B(n406), .Y(n493) );
  AO21_X0P5M_A12TR U768 ( .A0(n407), .A1(n406), .B0(n493), .Y(n448) );
  ADDF_X1M_A12TR U769 ( .A(b_s1[15]), .B(b_s1[16]), .CI(n408), .CO(n422), .S(
        n1335) );
  INV_X0P5B_A12TR U770 ( .A(b_s1[16]), .Y(n1086) );
  AOI22_X0P5M_A12TR U771 ( .A0(n1376), .A1(b_s1[15]), .B0(b_s1[17]), .B1(n1375), .Y(n409) );
  OAI211_X0P5M_A12TR U772 ( .A0(n1086), .A1(n1370), .B0(a_s1[2]), .C0(n409), 
        .Y(n411) );
  AOI22_X0P5M_A12TR U773 ( .A0(n1157), .A1(n1085), .B0(n1156), .B1(b_s1[17]), 
        .Y(n410) );
  AO21A1AI2_X0P5M_A12TR U774 ( .A0(n1085), .A1(n1141), .B0(n411), .C0(n410), 
        .Y(n412) );
  AOI21_X0P5M_A12TR U775 ( .A0(n1162), .A1(b_s1[16]), .B0(n412), .Y(n419) );
  XOR2_X0P5M_A12TR U776 ( .A(n420), .B(n419), .Y(n417) );
  CGENI_X1M_A12TR U777 ( .A(n415), .B(n414), .CI(n413), .CON(n418) );
  OAI21_X0P5M_A12TR U778 ( .A0(n417), .A1(n418), .B0(n1450), .Y(n416) );
  AOI21_X0P5M_A12TR U779 ( .A0(n417), .A1(n418), .B0(n416), .Y(
        \outreg_stage2/N20 ) );
  INV_X0P5B_A12TR U780 ( .A(n418), .Y(n421) );
  CGEN_X1M_A12TR U781 ( .A(n421), .B(n420), .CI(n419), .CO(n510) );
  ADDF_X1M_A12TR U782 ( .A(b_s1[16]), .B(b_s1[17]), .CI(n422), .CO(n503), .S(
        n1085) );
  INV_X0P5B_A12TR U783 ( .A(b_s1[17]), .Y(n1217) );
  AOI22_X0P5M_A12TR U784 ( .A0(n1376), .A1(b_s1[16]), .B0(b_s1[18]), .B1(n1375), .Y(n423) );
  OAI211_X0P5M_A12TR U785 ( .A0(n1217), .A1(n1370), .B0(a_s1[2]), .C0(n423), 
        .Y(n425) );
  AOI22_X0P5M_A12TR U786 ( .A0(n1157), .A1(n1214), .B0(n1156), .B1(b_s1[18]), 
        .Y(n424) );
  AO21A1AI2_X0P5M_A12TR U787 ( .A0(n1214), .A1(n1373), .B0(n425), .C0(n424), 
        .Y(n426) );
  AOI21_X0P5M_A12TR U788 ( .A0(n1162), .A1(b_s1[17]), .B0(n426), .Y(n509) );
  ADDF_X1M_A12TR U789 ( .A(n429), .B(n428), .CI(n427), .CO(n466), .S(n420) );
  OAI22_X0P5M_A12TR U790 ( .A0(n1168), .A1(n1235), .B0(n1167), .B1(n1237), .Y(
        n433) );
  AOI22_X0P5M_A12TR U791 ( .A0(n1301), .A1(n1233), .B0(n1302), .B1(b_s1[15]), 
        .Y(n430) );
  OAI211_X0P5M_A12TR U792 ( .A0(n1235), .A1(n1170), .B0(a_s1[5]), .C0(n430), 
        .Y(n431) );
  OAI222_X0P5M_A12TR U793 ( .A0(n431), .A1(n1299), .B0(n431), .B1(b_s1[13]), 
        .C0(n1173), .C1(n1098), .Y(n432) );
  AOI211_X0P5M_A12TR U794 ( .A0(n1178), .A1(n1233), .B0(n433), .C0(n432), .Y(
        n465) );
  ADDF_X1M_A12TR U795 ( .A(n436), .B(n435), .CI(n434), .CO(n473), .S(n427) );
  OAI22_X0P5M_A12TR U796 ( .A0(n971), .A1(n1184), .B0(n1025), .B1(n1182), .Y(
        n440) );
  AOI22_X0P5M_A12TR U797 ( .A0(n1359), .A1(n1267), .B0(n1362), .B1(b_s1[12]), 
        .Y(n437) );
  OAI211_X0P5M_A12TR U798 ( .A0(n971), .A1(n1187), .B0(a_s1[8]), .C0(n437), 
        .Y(n438) );
  OAI222_X0P5M_A12TR U799 ( .A0(n438), .A1(n1358), .B0(n438), .B1(b_s1[10]), 
        .C0(n1189), .C1(n892), .Y(n439) );
  AOI211_X0P5M_A12TR U800 ( .A0(n1194), .A1(n1267), .B0(n440), .C0(n439), .Y(
        n472) );
  ADDF_X1M_A12TR U801 ( .A(n443), .B(n442), .CI(n441), .CO(n480), .S(n434) );
  OAI22_X0P5M_A12TR U802 ( .A0(n782), .A1(n1200), .B0(n829), .B1(n1198), .Y(
        n447) );
  AOI22_X0P5M_A12TR U803 ( .A0(n1325), .A1(n1260), .B0(n1328), .B1(b_s1[9]), 
        .Y(n444) );
  OAI211_X0P5M_A12TR U804 ( .A0(n782), .A1(n1203), .B0(a_s1[11]), .C0(n444), 
        .Y(n445) );
  AOI211_X0P5M_A12TR U805 ( .A0(n1210), .A1(n1260), .B0(n447), .C0(n446), .Y(
        n479) );
  ADDF_X1M_A12TR U806 ( .A(n450), .B(n449), .CI(n448), .CO(n487), .S(n441) );
  INV_X0P5B_A12TR U807 ( .A(n1253), .Y(n612) );
  OAI22_X0P5M_A12TR U808 ( .A0(n614), .A1(n1216), .B0(n1215), .B1(n612), .Y(
        n454) );
  AOI22_X0P5M_A12TR U809 ( .A0(b_s1[4]), .A1(n1304), .B0(n1305), .B1(n1253), 
        .Y(n451) );
  OAI211_X0P5M_A12TR U810 ( .A0(n614), .A1(n883), .B0(a_s1[14]), .C0(n451), 
        .Y(n452) );
  AOI211_X0P5M_A12TR U811 ( .A0(b_s1[4]), .A1(n1226), .B0(n454), .C0(n453), 
        .Y(n486) );
  INV_X0P5B_A12TR U812 ( .A(n455), .Y(n1242) );
  OAI22_X0P5M_A12TR U813 ( .A0(n456), .A1(n1231), .B0(n458), .B1(n1232), .Y(
        n462) );
  INV_X0P5B_A12TR U814 ( .A(n1338), .Y(n1236) );
  AOI22_X0P5M_A12TR U815 ( .A0(n1243), .A1(n1334), .B0(b_s1[1]), .B1(n1336), 
        .Y(n457) );
  OAI211_X0P5M_A12TR U816 ( .A0(n458), .A1(n1236), .B0(a_s1[17]), .C0(n457), 
        .Y(n460) );
  INV_X0P5B_A12TR U817 ( .A(n459), .Y(n1238) );
  AOI211_X0P5M_A12TR U818 ( .A0(b_s1[1]), .A1(n1242), .B0(n462), .C0(n461), 
        .Y(n492) );
  INV_X0P5B_A12TR U819 ( .A(n551), .Y(n500) );
  NOR2_X0P5B_A12TR U820 ( .A(n1247), .B(n500), .Y(n556) );
  XOR3_X0P5M_A12TR U821 ( .A(n492), .B(n493), .C(n556), .Y(n485) );
  NOR2_X0P5B_A12TR U822 ( .A(reset), .B(n463), .Y(\outreg_stage2/N21 ) );
  ADDF_X1M_A12TR U823 ( .A(n466), .B(n465), .CI(n464), .CO(n515), .S(n508) );
  OAI22_X0P5M_A12TR U824 ( .A0(n1168), .A1(n1237), .B0(n1167), .B1(n1086), .Y(
        n470) );
  AOI22_X0P5M_A12TR U825 ( .A0(n1301), .A1(n1335), .B0(n1302), .B1(b_s1[16]), 
        .Y(n467) );
  OAI211_X0P5M_A12TR U826 ( .A0(n1237), .A1(n1170), .B0(a_s1[5]), .C0(n467), 
        .Y(n468) );
  OAI222_X0P5M_A12TR U827 ( .A0(n468), .A1(n1299), .B0(n468), .B1(b_s1[14]), 
        .C0(n1173), .C1(n1235), .Y(n469) );
  AOI211_X0P5M_A12TR U828 ( .A0(n1178), .A1(n1335), .B0(n470), .C0(n469), .Y(
        n514) );
  ADDF_X1M_A12TR U829 ( .A(n473), .B(n472), .CI(n471), .CO(n522), .S(n464) );
  OAI22_X0P5M_A12TR U830 ( .A0(n1025), .A1(n1184), .B0(n1098), .B1(n1182), .Y(
        n477) );
  AOI22_X0P5M_A12TR U831 ( .A0(n1359), .A1(n1312), .B0(n1362), .B1(b_s1[13]), 
        .Y(n474) );
  OAI211_X0P5M_A12TR U832 ( .A0(n1025), .A1(n1187), .B0(a_s1[8]), .C0(n474), 
        .Y(n475) );
  OAI222_X0P5M_A12TR U833 ( .A0(n475), .A1(n1358), .B0(n475), .B1(b_s1[11]), 
        .C0(n1189), .C1(n971), .Y(n476) );
  AOI211_X0P5M_A12TR U834 ( .A0(n1312), .A1(n1194), .B0(n477), .C0(n476), .Y(
        n521) );
  ADDF_X1M_A12TR U835 ( .A(n480), .B(n479), .CI(n478), .CO(n529), .S(n471) );
  OAI22_X0P5M_A12TR U836 ( .A0(n892), .A1(n1198), .B0(n829), .B1(n1200), .Y(
        n484) );
  AOI22_X0P5M_A12TR U837 ( .A0(n1325), .A1(n1332), .B0(n1328), .B1(b_s1[10]), 
        .Y(n481) );
  OAI211_X0P5M_A12TR U838 ( .A0(n829), .A1(n1203), .B0(a_s1[11]), .C0(n481), 
        .Y(n482) );
  AOI211_X0P5M_A12TR U839 ( .A0(n1332), .A1(n1210), .B0(n484), .C0(n483), .Y(
        n528) );
  ADDF_X1M_A12TR U840 ( .A(n487), .B(n486), .CI(n485), .CO(n536), .S(n478) );
  INV_X0P5B_A12TR U841 ( .A(n1378), .Y(n653) );
  OAI22_X0P5M_A12TR U842 ( .A0(n653), .A1(n1215), .B0(n655), .B1(n1216), .Y(
        n491) );
  AOI22_X0P5M_A12TR U843 ( .A0(b_s1[5]), .A1(n1304), .B0(n1378), .B1(n1305), 
        .Y(n488) );
  OAI211_X0P5M_A12TR U844 ( .A0(n655), .A1(n883), .B0(a_s1[14]), .C0(n488), 
        .Y(n489) );
  AOI211_X0P5M_A12TR U845 ( .A0(b_s1[5]), .A1(n1226), .B0(n491), .C0(n490), 
        .Y(n535) );
  OAI21B_X0P5M_A12TR U846 ( .A0(n556), .A1(n493), .B0N(n492), .Y(n543) );
  OAI22_X0P5M_A12TR U847 ( .A0(n496), .A1(n1232), .B0(n494), .B1(n1231), .Y(
        n499) );
  AOI22_X0P5M_A12TR U848 ( .A0(b_s1[2]), .A1(n1336), .B0(n1342), .B1(n1334), 
        .Y(n495) );
  OAI211_X0P5M_A12TR U849 ( .A0(n496), .A1(n1236), .B0(a_s1[17]), .C0(n495), 
        .Y(n497) );
  AOI211_X0P5M_A12TR U850 ( .A0(b_s1[2]), .A1(n1242), .B0(n499), .C0(n498), 
        .Y(n542) );
  NOR2_X0P5B_A12TR U851 ( .A(n550), .B(n500), .Y(n1311) );
  NOR2XB_X0P5M_A12TR U852 ( .BN(n550), .A(n500), .Y(n1309) );
  XOR2_X0P5M_A12TR U853 ( .A(a_s1[19]), .B(a_s1[18]), .Y(n552) );
  NOR2XB_X0P5M_A12TR U854 ( .BN(n552), .A(n551), .Y(n1310) );
  AOI222_X0P5M_A12TR U855 ( .A0(n1311), .A1(n1298), .B0(n1309), .B1(b_s1[1]), 
        .C0(n1310), .C1(b_s1[0]), .Y(n501) );
  INV_X0P5B_A12TR U856 ( .A(n501), .Y(n557) );
  NAND3_X0P5M_A12TR U857 ( .A(n556), .B(a_s1[20]), .C(n557), .Y(n502) );
  AO21A1AI2_X0P5M_A12TR U858 ( .A0(a_s1[20]), .A1(n556), .B0(n557), .C0(n502), 
        .Y(n541) );
  ADDF_X1M_A12TR U859 ( .A(b_s1[17]), .B(b_s1[18]), .CI(n503), .CO(n562), .S(
        n1214) );
  INV_X0P5B_A12TR U860 ( .A(b_s1[18]), .Y(n1221) );
  AOI22_X0P5M_A12TR U861 ( .A0(n1376), .A1(b_s1[17]), .B0(b_s1[19]), .B1(n1375), .Y(n504) );
  OAI211_X0P5M_A12TR U862 ( .A0(n1221), .A1(n1370), .B0(a_s1[2]), .C0(n504), 
        .Y(n506) );
  AOI22_X0P5M_A12TR U863 ( .A0(n1157), .A1(n1306), .B0(n1156), .B1(b_s1[19]), 
        .Y(n505) );
  AO21A1AI2_X0P5M_A12TR U864 ( .A0(n1306), .A1(n1141), .B0(n506), .C0(n505), 
        .Y(n507) );
  AOI21_X0P5M_A12TR U865 ( .A0(n1162), .A1(b_s1[18]), .B0(n507), .Y(n568) );
  ADDF_X1M_A12TR U866 ( .A(n510), .B(n509), .CI(n508), .CO(n567), .S(n463) );
  XNOR2_X0P5M_A12TR U867 ( .A(n568), .B(n567), .Y(n512) );
  OAI21_X0P5M_A12TR U868 ( .A0(n569), .A1(n512), .B0(n1450), .Y(n511) );
  AOI21_X0P5M_A12TR U869 ( .A0(n569), .A1(n512), .B0(n511), .Y(
        \outreg_stage2/N22 ) );
  ADDF_X1M_A12TR U870 ( .A(n515), .B(n514), .CI(n513), .CO(n583), .S(n569) );
  OAI22_X0P5M_A12TR U871 ( .A0(n1168), .A1(n1086), .B0(n1167), .B1(n1217), .Y(
        n519) );
  AOI22_X0P5M_A12TR U872 ( .A0(n1301), .A1(n1085), .B0(n1302), .B1(b_s1[17]), 
        .Y(n516) );
  OAI211_X0P5M_A12TR U873 ( .A0(n1086), .A1(n1170), .B0(a_s1[5]), .C0(n516), 
        .Y(n517) );
  OAI222_X0P5M_A12TR U874 ( .A0(n517), .A1(n1299), .B0(n517), .B1(b_s1[15]), 
        .C0(n1173), .C1(n1237), .Y(n518) );
  AOI211_X0P5M_A12TR U875 ( .A0(n1178), .A1(n1085), .B0(n519), .C0(n518), .Y(
        n582) );
  ADDF_X1M_A12TR U876 ( .A(n522), .B(n521), .CI(n520), .CO(n590), .S(n513) );
  OAI22_X0P5M_A12TR U877 ( .A0(n1098), .A1(n1184), .B0(n1235), .B1(n1182), .Y(
        n526) );
  AOI22_X0P5M_A12TR U878 ( .A0(n1359), .A1(n1096), .B0(n1362), .B1(b_s1[14]), 
        .Y(n523) );
  OAI211_X0P5M_A12TR U879 ( .A0(n1098), .A1(n1187), .B0(a_s1[8]), .C0(n523), 
        .Y(n524) );
  OAI222_X0P5M_A12TR U880 ( .A0(n524), .A1(n1358), .B0(n524), .B1(b_s1[12]), 
        .C0(n1189), .C1(n1025), .Y(n525) );
  AOI211_X0P5M_A12TR U881 ( .A0(n1194), .A1(n1096), .B0(n526), .C0(n525), .Y(
        n589) );
  ADDF_X1M_A12TR U882 ( .A(n529), .B(n528), .CI(n527), .CO(n597), .S(n520) );
  OAI22_X0P5M_A12TR U883 ( .A0(n971), .A1(n1198), .B0(n892), .B1(n1200), .Y(
        n533) );
  AOI22_X0P5M_A12TR U884 ( .A0(b_s1[11]), .A1(n1328), .B0(n1325), .B1(n1132), 
        .Y(n530) );
  OAI211_X0P5M_A12TR U885 ( .A0(n892), .A1(n1203), .B0(a_s1[11]), .C0(n530), 
        .Y(n531) );
  AOI211_X0P5M_A12TR U886 ( .A0(n1210), .A1(n1132), .B0(n533), .C0(n532), .Y(
        n596) );
  ADDF_X1M_A12TR U887 ( .A(n536), .B(n535), .CI(n534), .CO(n604), .S(n527) );
  INV_X0P5B_A12TR U888 ( .A(n1125), .Y(n707) );
  OAI22_X0P5M_A12TR U889 ( .A0(n709), .A1(n1216), .B0(n1215), .B1(n707), .Y(
        n540) );
  AOI22_X0P5M_A12TR U890 ( .A0(b_s1[6]), .A1(n1304), .B0(n1305), .B1(n1125), 
        .Y(n537) );
  OAI211_X0P5M_A12TR U891 ( .A0(n709), .A1(n883), .B0(a_s1[14]), .C0(n537), 
        .Y(n538) );
  AOI211_X0P5M_A12TR U892 ( .A0(b_s1[6]), .A1(n1226), .B0(n540), .C0(n539), 
        .Y(n603) );
  ADDF_X1M_A12TR U893 ( .A(n543), .B(n542), .CI(n541), .CO(n611), .S(n534) );
  OAI22_X0P5M_A12TR U894 ( .A0(n546), .A1(n1232), .B0(n544), .B1(n1231), .Y(
        n549) );
  AOI22_X0P5M_A12TR U895 ( .A0(b_s1[3]), .A1(n1336), .B0(n1118), .B1(n1334), 
        .Y(n545) );
  OAI211_X0P5M_A12TR U896 ( .A0(n546), .A1(n1236), .B0(a_s1[17]), .C0(n545), 
        .Y(n547) );
  AOI211_X0P5M_A12TR U897 ( .A0(b_s1[3]), .A1(n1242), .B0(n549), .C0(n548), 
        .Y(n610) );
  NOR3_X0P7M_A12TR U898 ( .A(n552), .B(n551), .C(n550), .Y(n1313) );
  AOI22_X0P5M_A12TR U899 ( .A0(b_s1[0]), .A1(n1313), .B0(n1109), .B1(n1311), 
        .Y(n555) );
  AOI22_X0P5M_A12TR U900 ( .A0(b_s1[1]), .A1(n1310), .B0(b_s1[2]), .B1(n1309), 
        .Y(n554) );
  INV_X0P5B_A12TR U901 ( .A(a_s1[20]), .Y(n1383) );
  NAND3_X0P5M_A12TR U902 ( .A(n554), .B(n555), .C(n1383), .Y(n553) );
  AO21A1AI2_X0P5M_A12TR U903 ( .A0(n555), .A1(n554), .B0(n1383), .C0(n553), 
        .Y(n561) );
  INV_X0P5B_A12TR U904 ( .A(n556), .Y(n559) );
  NOR2_X0P5B_A12TR U905 ( .A(n1383), .B(n557), .Y(n558) );
  NAND2_X0P5A_A12TR U906 ( .A(n559), .B(n558), .Y(n560) );
  NOR2_X0P5B_A12TR U907 ( .A(n561), .B(n560), .Y(n661) );
  AO21_X0P5M_A12TR U908 ( .A0(n561), .A1(n560), .B0(n661), .Y(n609) );
  ADDF_X1M_A12TR U909 ( .A(b_s1[18]), .B(b_s1[19]), .CI(n562), .CO(n576), .S(
        n1306) );
  INV_X0P5B_A12TR U910 ( .A(b_s1[19]), .Y(n1204) );
  AOI22_X0P5M_A12TR U911 ( .A0(n1376), .A1(b_s1[18]), .B0(b_s1[20]), .B1(n1375), .Y(n563) );
  OAI211_X0P5M_A12TR U912 ( .A0(n1204), .A1(n1370), .B0(a_s1[2]), .C0(n563), 
        .Y(n565) );
  AOI22_X0P5M_A12TR U913 ( .A0(n1157), .A1(n1081), .B0(n1156), .B1(b_s1[20]), 
        .Y(n564) );
  AO21A1AI2_X0P5M_A12TR U914 ( .A0(n1081), .A1(n1373), .B0(n565), .C0(n564), 
        .Y(n566) );
  AOI21_X0P5M_A12TR U915 ( .A0(n1162), .A1(b_s1[19]), .B0(n566), .Y(n573) );
  XOR2_X0P5M_A12TR U916 ( .A(n574), .B(n573), .Y(n571) );
  CGENI_X1M_A12TR U917 ( .A(n569), .B(n568), .CI(n567), .CON(n572) );
  OAI21_X0P5M_A12TR U918 ( .A0(n571), .A1(n572), .B0(n1450), .Y(n570) );
  AOI21_X0P5M_A12TR U919 ( .A0(n571), .A1(n572), .B0(n570), .Y(
        \outreg_stage2/N23 ) );
  INV_X0P5B_A12TR U920 ( .A(n572), .Y(n575) );
  CGEN_X1M_A12TR U921 ( .A(n575), .B(n574), .CI(n573), .CO(n673) );
  ADDF_X1M_A12TR U922 ( .A(b_s1[19]), .B(b_s1[20]), .CI(n576), .CO(n666), .S(
        n1081) );
  INV_X0P5B_A12TR U923 ( .A(b_s1[20]), .Y(n1202) );
  AOI22_X0P5M_A12TR U924 ( .A0(n1376), .A1(b_s1[19]), .B0(b_s1[21]), .B1(n1375), .Y(n577) );
  OAI211_X0P5M_A12TR U925 ( .A0(n1202), .A1(n1370), .B0(a_s1[2]), .C0(n577), 
        .Y(n579) );
  AOI22_X0P5M_A12TR U926 ( .A0(n1157), .A1(n1209), .B0(n1156), .B1(b_s1[21]), 
        .Y(n578) );
  AO21A1AI2_X0P5M_A12TR U927 ( .A0(n1209), .A1(n1141), .B0(n579), .C0(n578), 
        .Y(n580) );
  AOI21_X0P5M_A12TR U928 ( .A0(n1162), .A1(b_s1[20]), .B0(n580), .Y(n672) );
  ADDF_X1M_A12TR U929 ( .A(n583), .B(n582), .CI(n581), .CO(n624), .S(n574) );
  OAI22_X0P5M_A12TR U930 ( .A0(n1168), .A1(n1217), .B0(n1167), .B1(n1221), .Y(
        n587) );
  AOI22_X0P5M_A12TR U931 ( .A0(n1301), .A1(n1214), .B0(n1302), .B1(b_s1[18]), 
        .Y(n584) );
  OAI211_X0P5M_A12TR U932 ( .A0(n1217), .A1(n1170), .B0(a_s1[5]), .C0(n584), 
        .Y(n585) );
  OAI222_X0P5M_A12TR U933 ( .A0(n585), .A1(n1299), .B0(n585), .B1(b_s1[16]), 
        .C0(n1173), .C1(n1086), .Y(n586) );
  AOI211_X0P5M_A12TR U934 ( .A0(n1178), .A1(n1214), .B0(n587), .C0(n586), .Y(
        n623) );
  ADDF_X1M_A12TR U935 ( .A(n590), .B(n589), .CI(n588), .CO(n631), .S(n581) );
  OAI22_X0P5M_A12TR U936 ( .A0(n1235), .A1(n1184), .B0(n1237), .B1(n1182), .Y(
        n594) );
  AOI22_X0P5M_A12TR U937 ( .A0(n1359), .A1(n1233), .B0(n1362), .B1(b_s1[15]), 
        .Y(n591) );
  OAI211_X0P5M_A12TR U938 ( .A0(n1235), .A1(n1187), .B0(a_s1[8]), .C0(n591), 
        .Y(n592) );
  OAI222_X0P5M_A12TR U939 ( .A0(n592), .A1(n1358), .B0(n592), .B1(b_s1[13]), 
        .C0(n1189), .C1(n1098), .Y(n593) );
  AOI211_X0P5M_A12TR U940 ( .A0(n1194), .A1(n1233), .B0(n594), .C0(n593), .Y(
        n630) );
  ADDF_X1M_A12TR U941 ( .A(n597), .B(n596), .CI(n595), .CO(n638), .S(n588) );
  OAI22_X0P5M_A12TR U942 ( .A0(n971), .A1(n1200), .B0(n1025), .B1(n1198), .Y(
        n601) );
  AOI22_X0P5M_A12TR U943 ( .A0(b_s1[12]), .A1(n1328), .B0(n1325), .B1(n1267), 
        .Y(n598) );
  OAI211_X0P5M_A12TR U944 ( .A0(n1203), .A1(n971), .B0(a_s1[11]), .C0(n598), 
        .Y(n599) );
  AOI211_X0P5M_A12TR U945 ( .A0(n1210), .A1(n1267), .B0(n601), .C0(n600), .Y(
        n637) );
  ADDF_X1M_A12TR U946 ( .A(n604), .B(n603), .CI(n602), .CO(n645), .S(n595) );
  INV_X0P5B_A12TR U947 ( .A(n1260), .Y(n780) );
  OAI22_X0P5M_A12TR U948 ( .A0(n782), .A1(n1216), .B0(n1215), .B1(n780), .Y(
        n608) );
  AOI22_X0P5M_A12TR U949 ( .A0(b_s1[7]), .A1(n1304), .B0(n1305), .B1(n1260), 
        .Y(n605) );
  OAI211_X0P5M_A12TR U950 ( .A0(n782), .A1(n883), .B0(a_s1[14]), .C0(n605), 
        .Y(n606) );
  AOI211_X0P5M_A12TR U951 ( .A0(b_s1[7]), .A1(n1226), .B0(n608), .C0(n607), 
        .Y(n644) );
  ADDF_X1M_A12TR U952 ( .A(n611), .B(n610), .CI(n609), .CO(n652), .S(n602) );
  OAI22_X0P5M_A12TR U953 ( .A0(n614), .A1(n1232), .B0(n1231), .B1(n612), .Y(
        n617) );
  AOI22_X0P5M_A12TR U954 ( .A0(b_s1[4]), .A1(n1336), .B0(n1334), .B1(n1253), 
        .Y(n613) );
  OAI211_X0P5M_A12TR U955 ( .A0(n614), .A1(n1236), .B0(a_s1[17]), .C0(n613), 
        .Y(n615) );
  AOI211_X0P5M_A12TR U956 ( .A0(b_s1[4]), .A1(n1242), .B0(n617), .C0(n616), 
        .Y(n651) );
  INV_X0P5B_A12TR U957 ( .A(n715), .Y(n716) );
  NOR2_X0P5B_A12TR U958 ( .A(n1247), .B(n716), .Y(n662) );
  AOI22_X0P5M_A12TR U959 ( .A0(n1243), .A1(n1311), .B0(b_s1[1]), .B1(n1313), 
        .Y(n620) );
  AOI22_X0P5M_A12TR U960 ( .A0(b_s1[3]), .A1(n1309), .B0(b_s1[2]), .B1(n1310), 
        .Y(n619) );
  NAND3_X0P5M_A12TR U961 ( .A(n619), .B(n620), .C(a_s1[20]), .Y(n618) );
  AO21A1AI2_X0P5M_A12TR U962 ( .A0(n620), .A1(n619), .B0(a_s1[20]), .C0(n618), 
        .Y(n660) );
  XNOR3_X0P5M_A12TR U963 ( .A(n662), .B(n661), .C(n660), .Y(n650) );
  NOR2_X0P5B_A12TR U964 ( .A(reset), .B(n621), .Y(\outreg_stage2/N24 ) );
  ADDF_X1M_A12TR U965 ( .A(n624), .B(n623), .CI(n622), .CO(n678), .S(n671) );
  OAI22_X0P5M_A12TR U966 ( .A0(n1168), .A1(n1221), .B0(n1167), .B1(n1204), .Y(
        n628) );
  AOI22_X0P5M_A12TR U967 ( .A0(n1301), .A1(n1306), .B0(n1302), .B1(b_s1[19]), 
        .Y(n625) );
  OAI211_X0P5M_A12TR U968 ( .A0(n1221), .A1(n1170), .B0(a_s1[5]), .C0(n625), 
        .Y(n626) );
  OAI222_X0P5M_A12TR U969 ( .A0(n626), .A1(n1299), .B0(n626), .B1(b_s1[17]), 
        .C0(n1173), .C1(n1217), .Y(n627) );
  AOI211_X0P5M_A12TR U970 ( .A0(n1178), .A1(n1306), .B0(n628), .C0(n627), .Y(
        n677) );
  ADDF_X1M_A12TR U971 ( .A(n631), .B(n630), .CI(n629), .CO(n685), .S(n622) );
  OAI22_X0P5M_A12TR U972 ( .A0(n1237), .A1(n1184), .B0(n1086), .B1(n1182), .Y(
        n635) );
  AOI22_X0P5M_A12TR U973 ( .A0(n1359), .A1(n1335), .B0(n1362), .B1(b_s1[16]), 
        .Y(n632) );
  OAI211_X0P5M_A12TR U974 ( .A0(n1237), .A1(n1187), .B0(a_s1[8]), .C0(n632), 
        .Y(n633) );
  OAI222_X0P5M_A12TR U975 ( .A0(n633), .A1(n1358), .B0(n633), .B1(b_s1[14]), 
        .C0(n1189), .C1(n1235), .Y(n634) );
  AOI211_X0P5M_A12TR U976 ( .A0(n1335), .A1(n1194), .B0(n635), .C0(n634), .Y(
        n684) );
  ADDF_X1M_A12TR U977 ( .A(n638), .B(n637), .CI(n636), .CO(n692), .S(n629) );
  OAI22_X0P5M_A12TR U978 ( .A0(n1025), .A1(n1200), .B0(n1098), .B1(n1198), .Y(
        n642) );
  AOI22_X0P5M_A12TR U979 ( .A0(n1312), .A1(n1325), .B0(b_s1[13]), .B1(n1328), 
        .Y(n639) );
  OAI211_X0P5M_A12TR U980 ( .A0(n1203), .A1(n1025), .B0(a_s1[11]), .C0(n639), 
        .Y(n640) );
  AOI211_X0P5M_A12TR U981 ( .A0(n1312), .A1(n1210), .B0(n642), .C0(n641), .Y(
        n691) );
  ADDF_X1M_A12TR U982 ( .A(n645), .B(n644), .CI(n643), .CO(n699), .S(n636) );
  INV_X0P5B_A12TR U983 ( .A(n1332), .Y(n827) );
  OAI22_X0P5M_A12TR U984 ( .A0(n829), .A1(n1216), .B0(n827), .B1(n1215), .Y(
        n649) );
  AOI22_X0P5M_A12TR U985 ( .A0(n1305), .A1(n1332), .B0(n1304), .B1(b_s1[8]), 
        .Y(n646) );
  OAI211_X0P5M_A12TR U986 ( .A0(n829), .A1(n883), .B0(a_s1[14]), .C0(n646), 
        .Y(n647) );
  OAI222_X0P5M_A12TR U987 ( .A0(n647), .A1(n1307), .B0(n647), .B1(b_s1[10]), 
        .C0(n1222), .C1(n892), .Y(n648) );
  AOI211_X0P5M_A12TR U988 ( .A0(b_s1[8]), .A1(n1226), .B0(n649), .C0(n648), 
        .Y(n698) );
  ADDF_X1M_A12TR U989 ( .A(n652), .B(n651), .CI(n650), .CO(n706), .S(n643) );
  OAI22_X0P5M_A12TR U990 ( .A0(n653), .A1(n1231), .B0(n655), .B1(n1232), .Y(
        n658) );
  AOI22_X0P5M_A12TR U991 ( .A0(b_s1[5]), .A1(n1336), .B0(n1378), .B1(n1334), 
        .Y(n654) );
  OAI211_X0P5M_A12TR U992 ( .A0(n655), .A1(n1236), .B0(a_s1[17]), .C0(n654), 
        .Y(n656) );
  AOI211_X0P5M_A12TR U993 ( .A0(b_s1[5]), .A1(n1242), .B0(n658), .C0(n657), 
        .Y(n705) );
  NAND2_X0P5A_A12TR U994 ( .A(n662), .B(a_s1[23]), .Y(n659) );
  INV_X0P5B_A12TR U995 ( .A(a_s1[23]), .Y(n1424) );
  NOR2_X0P5B_A12TR U996 ( .A(n717), .B(n716), .Y(n1329) );
  XNOR2_X0P5M_A12TR U997 ( .A(a_s1[22]), .B(a_s1[21]), .Y(n718) );
  NOR2_X0P5B_A12TR U998 ( .A(n715), .B(n718), .Y(n1333) );
  AND2_X0P5M_A12TR U999 ( .A(n717), .B(n715), .Y(n1331) );
  AOI222_X0P5M_A12TR U1000 ( .A0(b_s1[1]), .A1(n1329), .B0(b_s1[0]), .B1(n1333), .C0(n1298), .C1(n1331), .Y(n713) );
  XNOR2_X0P5M_A12TR U1001 ( .A(n659), .B(n713), .Y(n726) );
  OAI21_X0P5M_A12TR U1002 ( .A0(n662), .A1(n661), .B0(n660), .Y(n725) );
  AOI22_X0P5M_A12TR U1003 ( .A0(b_s1[2]), .A1(n1313), .B0(n1342), .B1(n1311), 
        .Y(n665) );
  AOI22_X0P5M_A12TR U1004 ( .A0(b_s1[3]), .A1(n1310), .B0(b_s1[4]), .B1(n1309), 
        .Y(n664) );
  NAND3_X0P5M_A12TR U1005 ( .A(n664), .B(n665), .C(n1383), .Y(n663) );
  AO21A1AI2_X0P5M_A12TR U1006 ( .A0(n665), .A1(n664), .B0(n1383), .C0(n663), 
        .Y(n724) );
  ADDF_X1M_A12TR U1007 ( .A(b_s1[20]), .B(b_s1[21]), .CI(n666), .CO(n730), .S(
        n1209) );
  INV_X0P5B_A12TR U1008 ( .A(b_s1[21]), .Y(n1199) );
  AOI22_X0P5M_A12TR U1009 ( .A0(n1376), .A1(b_s1[20]), .B0(b_s1[22]), .B1(
        n1375), .Y(n667) );
  OAI211_X0P5M_A12TR U1010 ( .A0(n1199), .A1(n1370), .B0(a_s1[2]), .C0(n667), 
        .Y(n669) );
  AOI22_X0P5M_A12TR U1011 ( .A0(n1157), .A1(n1326), .B0(n1156), .B1(b_s1[22]), 
        .Y(n668) );
  AO21A1AI2_X0P5M_A12TR U1012 ( .A0(n1326), .A1(n1373), .B0(n669), .C0(n668), 
        .Y(n670) );
  AOI21_X0P5M_A12TR U1013 ( .A0(n1162), .A1(b_s1[21]), .B0(n670), .Y(n736) );
  ADDF_X1M_A12TR U1014 ( .A(n673), .B(n672), .CI(n671), .CO(n735), .S(n621) );
  XNOR2_X0P5M_A12TR U1015 ( .A(n736), .B(n735), .Y(n675) );
  OAI21_X0P5M_A12TR U1016 ( .A0(n737), .A1(n675), .B0(n1450), .Y(n674) );
  AOI21_X0P5M_A12TR U1017 ( .A0(n737), .A1(n675), .B0(n674), .Y(
        \outreg_stage2/N25 ) );
  ADDF_X1M_A12TR U1018 ( .A(n678), .B(n677), .CI(n676), .CO(n751), .S(n737) );
  OAI22_X0P5M_A12TR U1019 ( .A0(n1168), .A1(n1204), .B0(n1167), .B1(n1202), 
        .Y(n682) );
  AOI22_X0P5M_A12TR U1020 ( .A0(n1301), .A1(n1081), .B0(n1302), .B1(b_s1[20]), 
        .Y(n679) );
  OAI211_X0P5M_A12TR U1021 ( .A0(n1204), .A1(n1170), .B0(a_s1[5]), .C0(n679), 
        .Y(n680) );
  OAI222_X0P5M_A12TR U1022 ( .A0(n680), .A1(n1299), .B0(n680), .B1(b_s1[18]), 
        .C0(n1173), .C1(n1221), .Y(n681) );
  AOI211_X0P5M_A12TR U1023 ( .A0(n1178), .A1(n1081), .B0(n682), .C0(n681), .Y(
        n750) );
  ADDF_X1M_A12TR U1024 ( .A(n685), .B(n684), .CI(n683), .CO(n758), .S(n676) );
  OAI22_X0P5M_A12TR U1025 ( .A0(n1217), .A1(n1182), .B0(n1086), .B1(n1184), 
        .Y(n689) );
  AOI22_X0P5M_A12TR U1026 ( .A0(n1359), .A1(n1085), .B0(n1362), .B1(b_s1[17]), 
        .Y(n686) );
  OAI211_X0P5M_A12TR U1027 ( .A0(n1086), .A1(n1187), .B0(a_s1[8]), .C0(n686), 
        .Y(n687) );
  OAI222_X0P5M_A12TR U1028 ( .A0(n687), .A1(n1358), .B0(n687), .B1(b_s1[15]), 
        .C0(n1189), .C1(n1237), .Y(n688) );
  AOI211_X0P5M_A12TR U1029 ( .A0(n1194), .A1(n1085), .B0(n689), .C0(n688), .Y(
        n757) );
  ADDF_X1M_A12TR U1030 ( .A(n692), .B(n691), .CI(n690), .CO(n765), .S(n683) );
  OAI22_X0P5M_A12TR U1031 ( .A0(n1098), .A1(n1200), .B0(n1235), .B1(n1198), 
        .Y(n696) );
  AOI22_X0P5M_A12TR U1032 ( .A0(n1325), .A1(n1096), .B0(n1328), .B1(b_s1[14]), 
        .Y(n693) );
  OAI211_X0P5M_A12TR U1033 ( .A0(n1203), .A1(n1098), .B0(a_s1[11]), .C0(n693), 
        .Y(n694) );
  AOI211_X0P5M_A12TR U1034 ( .A0(n1210), .A1(n1096), .B0(n696), .C0(n695), .Y(
        n764) );
  ADDF_X1M_A12TR U1035 ( .A(n699), .B(n698), .CI(n697), .CO(n772), .S(n690) );
  INV_X0P5B_A12TR U1036 ( .A(n1132), .Y(n890) );
  OAI22_X0P5M_A12TR U1037 ( .A0(n892), .A1(n1216), .B0(n1215), .B1(n890), .Y(
        n703) );
  AOI22_X0P5M_A12TR U1038 ( .A0(n1305), .A1(n1132), .B0(n1304), .B1(b_s1[9]), 
        .Y(n700) );
  OAI211_X0P5M_A12TR U1039 ( .A0(n892), .A1(n883), .B0(a_s1[14]), .C0(n700), 
        .Y(n701) );
  OAI222_X0P5M_A12TR U1040 ( .A0(n701), .A1(n1307), .B0(n701), .B1(b_s1[11]), 
        .C0(n1222), .C1(n971), .Y(n702) );
  AOI211_X0P5M_A12TR U1041 ( .A0(b_s1[9]), .A1(n1226), .B0(n703), .C0(n702), 
        .Y(n771) );
  ADDF_X1M_A12TR U1042 ( .A(n706), .B(n705), .CI(n704), .CO(n779), .S(n697) );
  OAI22_X0P5M_A12TR U1043 ( .A0(n709), .A1(n1232), .B0(n1231), .B1(n707), .Y(
        n712) );
  AOI22_X0P5M_A12TR U1044 ( .A0(b_s1[6]), .A1(n1336), .B0(n1334), .B1(n1125), 
        .Y(n708) );
  OAI211_X0P5M_A12TR U1045 ( .A0(n709), .A1(n1236), .B0(a_s1[17]), .C0(n708), 
        .Y(n710) );
  AOI211_X0P5M_A12TR U1046 ( .A0(b_s1[6]), .A1(n1242), .B0(n712), .C0(n711), 
        .Y(n778) );
  INV_X0P5B_A12TR U1047 ( .A(n713), .Y(n714) );
  AOI211_X0P5M_A12TR U1048 ( .A0(b_s1[0]), .A1(n715), .B0(n1424), .C0(n714), 
        .Y(n723) );
  AND3_X0P5M_A12TR U1049 ( .A(n718), .B(n717), .C(n716), .Y(n1330) );
  AOI22_X0P5M_A12TR U1050 ( .A0(b_s1[2]), .A1(n1329), .B0(b_s1[0]), .B1(n1330), 
        .Y(n721) );
  AOI22_X0P5M_A12TR U1051 ( .A0(b_s1[1]), .A1(n1333), .B0(n1109), .B1(n1331), 
        .Y(n720) );
  NAND3_X0P5M_A12TR U1052 ( .A(n720), .B(n721), .C(a_s1[23]), .Y(n719) );
  AO21A1AI2_X0P5M_A12TR U1053 ( .A0(n721), .A1(n720), .B0(a_s1[23]), .C0(n719), 
        .Y(n722) );
  NAND2_X0P5A_A12TR U1054 ( .A(n723), .B(n722), .Y(n836) );
  OAI21_X0P5M_A12TR U1055 ( .A0(n723), .A1(n722), .B0(n836), .Y(n791) );
  ADDF_X1M_A12TR U1056 ( .A(n726), .B(n725), .CI(n724), .CO(n790), .S(n704) );
  AOI22_X0P5M_A12TR U1057 ( .A0(b_s1[3]), .A1(n1313), .B0(n1118), .B1(n1311), 
        .Y(n729) );
  AOI22_X0P5M_A12TR U1058 ( .A0(b_s1[4]), .A1(n1310), .B0(b_s1[5]), .B1(n1309), 
        .Y(n728) );
  NAND3_X0P5M_A12TR U1059 ( .A(n728), .B(n729), .C(n1383), .Y(n727) );
  AO21A1AI2_X0P5M_A12TR U1060 ( .A0(n729), .A1(n728), .B0(n1383), .C0(n727), 
        .Y(n789) );
  ADDF_X1M_A12TR U1061 ( .A(b_s1[21]), .B(b_s1[22]), .CI(n730), .CO(n744), .S(
        n1326) );
  INV_X0P5B_A12TR U1062 ( .A(b_s1[22]), .Y(n1188) );
  AOI22_X0P5M_A12TR U1063 ( .A0(n1376), .A1(b_s1[21]), .B0(b_s1[23]), .B1(
        n1375), .Y(n731) );
  OAI211_X0P5M_A12TR U1064 ( .A0(n1188), .A1(n1370), .B0(a_s1[2]), .C0(n731), 
        .Y(n733) );
  AOI22_X0P5M_A12TR U1065 ( .A0(n1157), .A1(n1073), .B0(n1156), .B1(b_s1[23]), 
        .Y(n732) );
  AO21A1AI2_X0P5M_A12TR U1066 ( .A0(n1073), .A1(n1141), .B0(n733), .C0(n732), 
        .Y(n734) );
  AOI21_X0P5M_A12TR U1067 ( .A0(n1162), .A1(b_s1[22]), .B0(n734), .Y(n741) );
  XOR2_X0P5M_A12TR U1068 ( .A(n742), .B(n741), .Y(n739) );
  CGENI_X1M_A12TR U1069 ( .A(n737), .B(n736), .CI(n735), .CON(n740) );
  OAI21_X0P5M_A12TR U1070 ( .A0(n739), .A1(n740), .B0(n1450), .Y(n738) );
  AOI21_X0P5M_A12TR U1071 ( .A0(n739), .A1(n740), .B0(n738), .Y(
        \outreg_stage2/N26 ) );
  INV_X0P5B_A12TR U1072 ( .A(n740), .Y(n743) );
  CGEN_X1M_A12TR U1073 ( .A(n743), .B(n742), .CI(n741), .CO(n855) );
  ADDF_X1M_A12TR U1074 ( .A(b_s1[22]), .B(b_s1[23]), .CI(n744), .CO(n848), .S(
        n1073) );
  INV_X0P5B_A12TR U1075 ( .A(b_s1[23]), .Y(n1186) );
  AOI22_X0P5M_A12TR U1076 ( .A0(n1376), .A1(b_s1[22]), .B0(b_s1[24]), .B1(
        n1375), .Y(n745) );
  OAI211_X0P5M_A12TR U1077 ( .A0(n1186), .A1(n1370), .B0(a_s1[2]), .C0(n745), 
        .Y(n747) );
  AOI22_X0P5M_A12TR U1078 ( .A0(n1157), .A1(n1193), .B0(n1156), .B1(b_s1[24]), 
        .Y(n746) );
  AO21A1AI2_X0P5M_A12TR U1079 ( .A0(n1193), .A1(n1373), .B0(n747), .C0(n746), 
        .Y(n748) );
  AOI21_X0P5M_A12TR U1080 ( .A0(n1162), .A1(b_s1[23]), .B0(n748), .Y(n854) );
  ADDF_X1M_A12TR U1081 ( .A(n751), .B(n750), .CI(n749), .CO(n798), .S(n742) );
  OAI22_X0P5M_A12TR U1082 ( .A0(n1168), .A1(n1202), .B0(n1167), .B1(n1199), 
        .Y(n755) );
  AOI22_X0P5M_A12TR U1083 ( .A0(n1301), .A1(n1209), .B0(n1302), .B1(b_s1[21]), 
        .Y(n752) );
  OAI211_X0P5M_A12TR U1084 ( .A0(n1202), .A1(n1170), .B0(a_s1[5]), .C0(n752), 
        .Y(n753) );
  OAI222_X0P5M_A12TR U1085 ( .A0(n753), .A1(n1299), .B0(n753), .B1(b_s1[19]), 
        .C0(n1173), .C1(n1204), .Y(n754) );
  AOI211_X0P5M_A12TR U1086 ( .A0(n1178), .A1(n1209), .B0(n755), .C0(n754), .Y(
        n797) );
  ADDF_X1M_A12TR U1087 ( .A(n758), .B(n757), .CI(n756), .CO(n805), .S(n749) );
  OAI22_X0P5M_A12TR U1088 ( .A0(n1217), .A1(n1184), .B0(n1221), .B1(n1182), 
        .Y(n762) );
  AOI22_X0P5M_A12TR U1089 ( .A0(n1359), .A1(n1214), .B0(n1362), .B1(b_s1[18]), 
        .Y(n759) );
  OAI211_X0P5M_A12TR U1090 ( .A0(n1217), .A1(n1187), .B0(a_s1[8]), .C0(n759), 
        .Y(n760) );
  OAI222_X0P5M_A12TR U1091 ( .A0(n760), .A1(n1358), .B0(n760), .B1(b_s1[16]), 
        .C0(n1189), .C1(n1086), .Y(n761) );
  AOI211_X0P5M_A12TR U1092 ( .A0(n1194), .A1(n1214), .B0(n762), .C0(n761), .Y(
        n804) );
  ADDF_X1M_A12TR U1093 ( .A(n765), .B(n764), .CI(n763), .CO(n812), .S(n756) );
  OAI22_X0P5M_A12TR U1094 ( .A0(n1235), .A1(n1200), .B0(n1237), .B1(n1198), 
        .Y(n769) );
  AOI22_X0P5M_A12TR U1095 ( .A0(n1325), .A1(n1233), .B0(n1328), .B1(b_s1[15]), 
        .Y(n766) );
  OAI211_X0P5M_A12TR U1096 ( .A0(n1235), .A1(n1203), .B0(a_s1[11]), .C0(n766), 
        .Y(n767) );
  AOI211_X0P5M_A12TR U1097 ( .A0(n1210), .A1(n1233), .B0(n769), .C0(n768), .Y(
        n811) );
  ADDF_X1M_A12TR U1098 ( .A(n772), .B(n771), .CI(n770), .CO(n819), .S(n763) );
  INV_X0P5B_A12TR U1099 ( .A(n1267), .Y(n969) );
  OAI22_X0P5M_A12TR U1100 ( .A0(n971), .A1(n1216), .B0(n1215), .B1(n969), .Y(
        n776) );
  AOI22_X0P5M_A12TR U1101 ( .A0(n1305), .A1(n1267), .B0(n1304), .B1(b_s1[10]), 
        .Y(n773) );
  OAI211_X0P5M_A12TR U1102 ( .A0(n971), .A1(n883), .B0(a_s1[14]), .C0(n773), 
        .Y(n774) );
  OAI222_X0P5M_A12TR U1103 ( .A0(n774), .A1(n1307), .B0(n774), .B1(b_s1[12]), 
        .C0(n1222), .C1(n1025), .Y(n775) );
  AOI211_X0P5M_A12TR U1104 ( .A0(b_s1[10]), .A1(n1226), .B0(n776), .C0(n775), 
        .Y(n818) );
  ADDF_X1M_A12TR U1105 ( .A(n779), .B(n778), .CI(n777), .CO(n826), .S(n770) );
  OAI22_X0P5M_A12TR U1106 ( .A0(n782), .A1(n1232), .B0(n1231), .B1(n780), .Y(
        n785) );
  AOI22_X0P5M_A12TR U1107 ( .A0(b_s1[7]), .A1(n1336), .B0(n1334), .B1(n1260), 
        .Y(n781) );
  OAI211_X0P5M_A12TR U1108 ( .A0(n1236), .A1(n782), .B0(a_s1[17]), .C0(n781), 
        .Y(n783) );
  AOI211_X0P5M_A12TR U1109 ( .A0(b_s1[7]), .A1(n1242), .B0(n785), .C0(n784), 
        .Y(n825) );
  INV_X0P5B_A12TR U1110 ( .A(n898), .Y(n900) );
  NOR2_X0P5B_A12TR U1111 ( .A(n1247), .B(n900), .Y(n837) );
  AOI22_X0P5M_A12TR U1112 ( .A0(b_s1[1]), .A1(n1330), .B0(b_s1[3]), .B1(n1329), 
        .Y(n788) );
  AOI22_X0P5M_A12TR U1113 ( .A0(n1243), .A1(n1331), .B0(b_s1[2]), .B1(n1333), 
        .Y(n787) );
  NAND3_X0P5M_A12TR U1114 ( .A(n787), .B(n788), .C(n1424), .Y(n786) );
  AO21A1AI2_X0P5M_A12TR U1115 ( .A0(n788), .A1(n787), .B0(n1424), .C0(n786), 
        .Y(n835) );
  XNOR3_X0P5M_A12TR U1116 ( .A(n837), .B(n835), .C(n836), .Y(n844) );
  ADDF_X1M_A12TR U1117 ( .A(n791), .B(n790), .CI(n789), .CO(n843), .S(n777) );
  AOI22_X0P5M_A12TR U1118 ( .A0(b_s1[4]), .A1(n1313), .B0(n1311), .B1(n1253), 
        .Y(n794) );
  AOI22_X0P5M_A12TR U1119 ( .A0(b_s1[5]), .A1(n1310), .B0(b_s1[6]), .B1(n1309), 
        .Y(n793) );
  NAND3_X0P5M_A12TR U1120 ( .A(n793), .B(n794), .C(n1383), .Y(n792) );
  AO21A1AI2_X0P5M_A12TR U1121 ( .A0(n794), .A1(n793), .B0(n1383), .C0(n792), 
        .Y(n842) );
  NOR2_X0P5B_A12TR U1122 ( .A(reset), .B(n795), .Y(\outreg_stage2/N27 ) );
  ADDF_X1M_A12TR U1123 ( .A(n798), .B(n797), .CI(n796), .CO(n860), .S(n853) );
  OAI22_X0P5M_A12TR U1124 ( .A0(n1168), .A1(n1199), .B0(n1167), .B1(n1188), 
        .Y(n802) );
  AOI22_X0P5M_A12TR U1125 ( .A0(n1301), .A1(n1326), .B0(n1302), .B1(b_s1[22]), 
        .Y(n799) );
  OAI211_X0P5M_A12TR U1126 ( .A0(n1199), .A1(n1170), .B0(a_s1[5]), .C0(n799), 
        .Y(n800) );
  OAI222_X0P5M_A12TR U1127 ( .A0(n800), .A1(n1299), .B0(n800), .B1(b_s1[20]), 
        .C0(n1173), .C1(n1202), .Y(n801) );
  AOI211_X0P5M_A12TR U1128 ( .A0(n1178), .A1(n1326), .B0(n802), .C0(n801), .Y(
        n859) );
  ADDF_X1M_A12TR U1129 ( .A(n805), .B(n804), .CI(n803), .CO(n867), .S(n796) );
  OAI22_X0P5M_A12TR U1130 ( .A0(n1221), .A1(n1184), .B0(n1204), .B1(n1182), 
        .Y(n809) );
  AOI22_X0P5M_A12TR U1131 ( .A0(n1359), .A1(n1306), .B0(n1362), .B1(b_s1[19]), 
        .Y(n806) );
  OAI211_X0P5M_A12TR U1132 ( .A0(n1221), .A1(n1187), .B0(a_s1[8]), .C0(n806), 
        .Y(n807) );
  OAI222_X0P5M_A12TR U1133 ( .A0(n807), .A1(n1358), .B0(n807), .B1(b_s1[17]), 
        .C0(n1189), .C1(n1217), .Y(n808) );
  AOI211_X0P5M_A12TR U1134 ( .A0(n1306), .A1(n1194), .B0(n809), .C0(n808), .Y(
        n866) );
  ADDF_X1M_A12TR U1135 ( .A(n812), .B(n811), .CI(n810), .CO(n874), .S(n803) );
  OAI22_X0P5M_A12TR U1136 ( .A0(n1237), .A1(n1200), .B0(n1086), .B1(n1198), 
        .Y(n816) );
  AOI22_X0P5M_A12TR U1137 ( .A0(n1325), .A1(n1335), .B0(n1328), .B1(b_s1[16]), 
        .Y(n813) );
  OAI211_X0P5M_A12TR U1138 ( .A0(n1237), .A1(n1203), .B0(a_s1[11]), .C0(n813), 
        .Y(n814) );
  AOI211_X0P5M_A12TR U1139 ( .A0(n1335), .A1(n1210), .B0(n816), .C0(n815), .Y(
        n873) );
  ADDF_X1M_A12TR U1140 ( .A(n819), .B(n818), .CI(n817), .CO(n881), .S(n810) );
  INV_X0P5B_A12TR U1141 ( .A(n1312), .Y(n1023) );
  OAI22_X0P5M_A12TR U1142 ( .A0(n1023), .A1(n1215), .B0(n1025), .B1(n1216), 
        .Y(n823) );
  AOI22_X0P5M_A12TR U1143 ( .A0(n1305), .A1(n1312), .B0(n1304), .B1(b_s1[11]), 
        .Y(n820) );
  OAI211_X0P5M_A12TR U1144 ( .A0(n1025), .A1(n883), .B0(a_s1[14]), .C0(n820), 
        .Y(n821) );
  OAI222_X0P5M_A12TR U1145 ( .A0(n821), .A1(n1307), .B0(n821), .B1(b_s1[13]), 
        .C0(n1222), .C1(n1098), .Y(n822) );
  AOI211_X0P5M_A12TR U1146 ( .A0(b_s1[11]), .A1(n1226), .B0(n823), .C0(n822), 
        .Y(n880) );
  ADDF_X1M_A12TR U1147 ( .A(n826), .B(n825), .CI(n824), .CO(n889), .S(n817) );
  OAI22_X0P5M_A12TR U1148 ( .A0(n829), .A1(n1232), .B0(n827), .B1(n1231), .Y(
        n832) );
  AOI22_X0P5M_A12TR U1149 ( .A0(b_s1[8]), .A1(n1336), .B0(n1332), .B1(n1334), 
        .Y(n828) );
  OAI211_X0P5M_A12TR U1150 ( .A0(n1236), .A1(n829), .B0(a_s1[17]), .C0(n828), 
        .Y(n830) );
  AOI211_X0P5M_A12TR U1151 ( .A0(b_s1[8]), .A1(n1242), .B0(n832), .C0(n831), 
        .Y(n888) );
  NAND2_X0P5A_A12TR U1152 ( .A(n837), .B(a_s1[26]), .Y(n834) );
  INV_X0P5B_A12TR U1153 ( .A(n833), .Y(n899) );
  NOR2_X0P5B_A12TR U1154 ( .A(n899), .B(n900), .Y(n1380) );
  XNOR2_X0P5M_A12TR U1155 ( .A(a_s1[25]), .B(a_s1[24]), .Y(n901) );
  NOR2_X0P5B_A12TR U1156 ( .A(n898), .B(n901), .Y(n1381) );
  NOR2_X0P5B_A12TR U1157 ( .A(n833), .B(n900), .Y(n1377) );
  AOI222_X0P5M_A12TR U1158 ( .A0(b_s1[1]), .A1(n1380), .B0(b_s1[0]), .B1(n1381), .C0(n1298), .C1(n1377), .Y(n896) );
  XNOR2_X0P5M_A12TR U1159 ( .A(n834), .B(n896), .Y(n909) );
  AOI2XB1_X0P5M_A12TR U1160 ( .A1N(n837), .A0(n836), .B0(n835), .Y(n838) );
  INV_X0P5B_A12TR U1161 ( .A(n838), .Y(n908) );
  AOI22_X0P5M_A12TR U1162 ( .A0(b_s1[2]), .A1(n1330), .B0(b_s1[4]), .B1(n1329), 
        .Y(n841) );
  AOI22_X0P5M_A12TR U1163 ( .A0(b_s1[3]), .A1(n1333), .B0(n1342), .B1(n1331), 
        .Y(n840) );
  NAND3_X0P5M_A12TR U1164 ( .A(n840), .B(n841), .C(n1424), .Y(n839) );
  AO21A1AI2_X0P5M_A12TR U1165 ( .A0(n841), .A1(n840), .B0(n1424), .C0(n839), 
        .Y(n907) );
  ADDF_X1M_A12TR U1166 ( .A(n844), .B(n843), .CI(n842), .CO(n914), .S(n824) );
  AOI22_X0P5M_A12TR U1167 ( .A0(b_s1[5]), .A1(n1313), .B0(n1378), .B1(n1311), 
        .Y(n847) );
  AOI22_X0P5M_A12TR U1168 ( .A0(b_s1[6]), .A1(n1310), .B0(b_s1[7]), .B1(n1309), 
        .Y(n846) );
  NAND3_X0P5M_A12TR U1169 ( .A(n846), .B(n847), .C(n1383), .Y(n845) );
  AO21A1AI2_X0P5M_A12TR U1170 ( .A0(n847), .A1(n846), .B0(n1383), .C0(n845), 
        .Y(n913) );
  ADDF_X1M_A12TR U1171 ( .A(b_s1[23]), .B(b_s1[24]), .CI(n848), .CO(n919), .S(
        n1193) );
  INV_X0P5B_A12TR U1172 ( .A(b_s1[24]), .Y(n1183) );
  AOI22_X0P5M_A12TR U1173 ( .A0(n1376), .A1(b_s1[23]), .B0(b_s1[25]), .B1(
        n1375), .Y(n849) );
  OAI211_X0P5M_A12TR U1174 ( .A0(n1183), .A1(n1370), .B0(a_s1[2]), .C0(n849), 
        .Y(n851) );
  AOI22_X0P5M_A12TR U1175 ( .A0(n1157), .A1(n1360), .B0(n1156), .B1(b_s1[25]), 
        .Y(n850) );
  AO21A1AI2_X0P5M_A12TR U1176 ( .A0(n1360), .A1(n1141), .B0(n851), .C0(n850), 
        .Y(n852) );
  AOI21_X0P5M_A12TR U1177 ( .A0(n1162), .A1(b_s1[24]), .B0(n852), .Y(n925) );
  ADDF_X1M_A12TR U1178 ( .A(n855), .B(n854), .CI(n853), .CO(n924), .S(n795) );
  XNOR2_X0P5M_A12TR U1179 ( .A(n925), .B(n924), .Y(n857) );
  OAI21_X0P5M_A12TR U1180 ( .A0(n926), .A1(n857), .B0(n1450), .Y(n856) );
  AOI21_X0P5M_A12TR U1181 ( .A0(n926), .A1(n857), .B0(n856), .Y(
        \outreg_stage2/N28 ) );
  ADDF_X1M_A12TR U1182 ( .A(n860), .B(n859), .CI(n858), .CO(n940), .S(n926) );
  OAI22_X0P5M_A12TR U1183 ( .A0(n1168), .A1(n1188), .B0(n1167), .B1(n1186), 
        .Y(n864) );
  AOI22_X0P5M_A12TR U1184 ( .A0(n1301), .A1(n1073), .B0(n1302), .B1(b_s1[23]), 
        .Y(n861) );
  OAI211_X0P5M_A12TR U1185 ( .A0(n1188), .A1(n1170), .B0(a_s1[5]), .C0(n861), 
        .Y(n862) );
  OAI222_X0P5M_A12TR U1186 ( .A0(n862), .A1(n1299), .B0(n862), .B1(b_s1[21]), 
        .C0(n1173), .C1(n1199), .Y(n863) );
  AOI211_X0P5M_A12TR U1187 ( .A0(n1178), .A1(n1073), .B0(n864), .C0(n863), .Y(
        n939) );
  ADDF_X1M_A12TR U1188 ( .A(n867), .B(n866), .CI(n865), .CO(n947), .S(n858) );
  OAI22_X0P5M_A12TR U1189 ( .A0(n1204), .A1(n1184), .B0(n1202), .B1(n1182), 
        .Y(n871) );
  AOI22_X0P5M_A12TR U1190 ( .A0(n1359), .A1(n1081), .B0(n1362), .B1(b_s1[20]), 
        .Y(n868) );
  OAI211_X0P5M_A12TR U1191 ( .A0(n1204), .A1(n1187), .B0(a_s1[8]), .C0(n868), 
        .Y(n869) );
  OAI222_X0P5M_A12TR U1192 ( .A0(n869), .A1(n1358), .B0(n869), .B1(b_s1[18]), 
        .C0(n1189), .C1(n1221), .Y(n870) );
  AOI211_X0P5M_A12TR U1193 ( .A0(n1194), .A1(n1081), .B0(n871), .C0(n870), .Y(
        n946) );
  ADDF_X1M_A12TR U1194 ( .A(n874), .B(n873), .CI(n872), .CO(n954), .S(n865) );
  OAI22_X0P5M_A12TR U1195 ( .A0(n1217), .A1(n1198), .B0(n1086), .B1(n1200), 
        .Y(n878) );
  AOI22_X0P5M_A12TR U1196 ( .A0(b_s1[17]), .A1(n1328), .B0(n1325), .B1(n1085), 
        .Y(n875) );
  OAI211_X0P5M_A12TR U1197 ( .A0(n1086), .A1(n1203), .B0(a_s1[11]), .C0(n875), 
        .Y(n876) );
  AOI211_X0P5M_A12TR U1198 ( .A0(n1210), .A1(n1085), .B0(n878), .C0(n877), .Y(
        n953) );
  ADDF_X1M_A12TR U1199 ( .A(n881), .B(n880), .CI(n879), .CO(n961), .S(n872) );
  INV_X0P5B_A12TR U1200 ( .A(n1096), .Y(n1095) );
  OAI22_X0P5M_A12TR U1201 ( .A0(n1098), .A1(n1216), .B0(n1215), .B1(n1095), 
        .Y(n886) );
  AOI22_X0P5M_A12TR U1202 ( .A0(n1305), .A1(n1096), .B0(n1304), .B1(b_s1[12]), 
        .Y(n882) );
  OAI211_X0P5M_A12TR U1203 ( .A0(n1098), .A1(n883), .B0(a_s1[14]), .C0(n882), 
        .Y(n884) );
  OAI222_X0P5M_A12TR U1204 ( .A0(n884), .A1(n1307), .B0(n884), .B1(b_s1[14]), 
        .C0(n1222), .C1(n1235), .Y(n885) );
  AOI211_X0P5M_A12TR U1205 ( .A0(b_s1[12]), .A1(n1226), .B0(n886), .C0(n885), 
        .Y(n960) );
  ADDF_X1M_A12TR U1206 ( .A(n889), .B(n888), .CI(n887), .CO(n968), .S(n879) );
  OAI22_X0P5M_A12TR U1207 ( .A0(n892), .A1(n1232), .B0(n1231), .B1(n890), .Y(
        n895) );
  AOI22_X0P5M_A12TR U1208 ( .A0(b_s1[9]), .A1(n1336), .B0(n1334), .B1(n1132), 
        .Y(n891) );
  OAI211_X0P5M_A12TR U1209 ( .A0(n1236), .A1(n892), .B0(a_s1[17]), .C0(n891), 
        .Y(n893) );
  AOI211_X0P5M_A12TR U1210 ( .A0(b_s1[9]), .A1(n1242), .B0(n895), .C0(n894), 
        .Y(n967) );
  NAND2_X0P5A_A12TR U1211 ( .A(a_s1[26]), .B(n896), .Y(n897) );
  AOI21_X0P5M_A12TR U1212 ( .A0(n898), .A1(b_s1[0]), .B0(n897), .Y(n906) );
  AND3_X0P5M_A12TR U1213 ( .A(n901), .B(n900), .C(n899), .Y(n1379) );
  AOI22_X0P5M_A12TR U1214 ( .A0(b_s1[0]), .A1(n1379), .B0(n1109), .B1(n1377), 
        .Y(n904) );
  AOI22_X0P5M_A12TR U1215 ( .A0(b_s1[1]), .A1(n1381), .B0(b_s1[2]), .B1(n1380), 
        .Y(n903) );
  NAND3_X0P5M_A12TR U1216 ( .A(n903), .B(n904), .C(a_s1[26]), .Y(n902) );
  AO21A1AI2_X0P5M_A12TR U1217 ( .A0(n904), .A1(n903), .B0(a_s1[26]), .C0(n902), 
        .Y(n905) );
  NAND2_X0P5A_A12TR U1218 ( .A(n906), .B(n905), .Y(n1032) );
  OAI21_X0P5M_A12TR U1219 ( .A0(n906), .A1(n905), .B0(n1032), .Y(n980) );
  ADDF_X1M_A12TR U1220 ( .A(n909), .B(n908), .CI(n907), .CO(n979), .S(n915) );
  AOI22_X0P5M_A12TR U1221 ( .A0(b_s1[3]), .A1(n1330), .B0(b_s1[5]), .B1(n1329), 
        .Y(n912) );
  AOI22_X0P5M_A12TR U1222 ( .A0(b_s1[4]), .A1(n1333), .B0(n1118), .B1(n1331), 
        .Y(n911) );
  NAND3_X0P5M_A12TR U1223 ( .A(n911), .B(n912), .C(n1424), .Y(n910) );
  AO21A1AI2_X0P5M_A12TR U1224 ( .A0(n912), .A1(n911), .B0(n1424), .C0(n910), 
        .Y(n978) );
  ADDF_X1M_A12TR U1225 ( .A(n915), .B(n914), .CI(n913), .CO(n985), .S(n887) );
  AOI22_X0P5M_A12TR U1226 ( .A0(b_s1[6]), .A1(n1313), .B0(n1311), .B1(n1125), 
        .Y(n918) );
  AOI22_X0P5M_A12TR U1227 ( .A0(b_s1[7]), .A1(n1310), .B0(n1309), .B1(b_s1[8]), 
        .Y(n917) );
  NAND3_X0P5M_A12TR U1228 ( .A(n917), .B(n918), .C(n1383), .Y(n916) );
  AO21A1AI2_X0P5M_A12TR U1229 ( .A0(n918), .A1(n917), .B0(n1383), .C0(n916), 
        .Y(n984) );
  ADDF_X1M_A12TR U1230 ( .A(b_s1[24]), .B(b_s1[25]), .CI(n919), .CO(n933), .S(
        n1360) );
  INV_X0P5B_A12TR U1231 ( .A(b_s1[25]), .Y(n1172) );
  AOI22_X0P5M_A12TR U1232 ( .A0(n1376), .A1(b_s1[24]), .B0(b_s1[26]), .B1(
        n1375), .Y(n920) );
  OAI211_X0P5M_A12TR U1233 ( .A0(n1172), .A1(n1370), .B0(a_s1[2]), .C0(n920), 
        .Y(n922) );
  AOI22_X0P5M_A12TR U1234 ( .A0(n1157), .A1(n1065), .B0(n1156), .B1(b_s1[26]), 
        .Y(n921) );
  AO21A1AI2_X0P5M_A12TR U1235 ( .A0(n1065), .A1(n1373), .B0(n922), .C0(n921), 
        .Y(n923) );
  AOI21_X0P5M_A12TR U1236 ( .A0(n1162), .A1(b_s1[25]), .B0(n923), .Y(n930) );
  XOR2_X0P5M_A12TR U1237 ( .A(n931), .B(n930), .Y(n928) );
  CGENI_X1M_A12TR U1238 ( .A(n926), .B(n925), .CI(n924), .CON(n929) );
  OAI21_X0P5M_A12TR U1239 ( .A0(n928), .A1(n929), .B0(n1450), .Y(n927) );
  AOI21_X0P5M_A12TR U1240 ( .A0(n928), .A1(n929), .B0(n927), .Y(
        \outreg_stage2/N29 ) );
  INV_X0P5B_A12TR U1241 ( .A(n929), .Y(n932) );
  CGEN_X1M_A12TR U1242 ( .A(n932), .B(n931), .CI(n930), .CO(n1055) );
  ADDF_X1M_A12TR U1243 ( .A(b_s1[25]), .B(b_s1[26]), .CI(n933), .CO(n1048), 
        .S(n1065) );
  INV_X0P5B_A12TR U1244 ( .A(b_s1[26]), .Y(n1171) );
  AOI22_X0P5M_A12TR U1245 ( .A0(n1376), .A1(b_s1[25]), .B0(b_s1[27]), .B1(
        n1375), .Y(n934) );
  OAI211_X0P5M_A12TR U1246 ( .A0(n1171), .A1(n1370), .B0(a_s1[2]), .C0(n934), 
        .Y(n936) );
  AOI22_X0P5M_A12TR U1247 ( .A0(n1157), .A1(n1177), .B0(n1156), .B1(b_s1[27]), 
        .Y(n935) );
  AO21A1AI2_X0P5M_A12TR U1248 ( .A0(n1177), .A1(n1141), .B0(n936), .C0(n935), 
        .Y(n937) );
  AOI21_X0P5M_A12TR U1249 ( .A0(n1162), .A1(b_s1[26]), .B0(n937), .Y(n1054) );
  ADDF_X1M_A12TR U1250 ( .A(n940), .B(n939), .CI(n938), .CO(n993), .S(n931) );
  OAI22_X0P5M_A12TR U1251 ( .A0(n1168), .A1(n1186), .B0(n1167), .B1(n1183), 
        .Y(n944) );
  AOI22_X0P5M_A12TR U1252 ( .A0(n1301), .A1(n1193), .B0(n1302), .B1(b_s1[24]), 
        .Y(n941) );
  OAI211_X0P5M_A12TR U1253 ( .A0(n1186), .A1(n1170), .B0(a_s1[5]), .C0(n941), 
        .Y(n942) );
  OAI222_X0P5M_A12TR U1254 ( .A0(n942), .A1(n1299), .B0(n942), .B1(b_s1[22]), 
        .C0(n1173), .C1(n1188), .Y(n943) );
  AOI211_X0P5M_A12TR U1255 ( .A0(n1178), .A1(n1193), .B0(n944), .C0(n943), .Y(
        n992) );
  ADDF_X1M_A12TR U1256 ( .A(n947), .B(n946), .CI(n945), .CO(n1000), .S(n938)
         );
  OAI22_X0P5M_A12TR U1257 ( .A0(n1202), .A1(n1184), .B0(n1199), .B1(n1182), 
        .Y(n951) );
  AOI22_X0P5M_A12TR U1258 ( .A0(n1359), .A1(n1209), .B0(n1362), .B1(b_s1[21]), 
        .Y(n948) );
  OAI211_X0P5M_A12TR U1259 ( .A0(n1202), .A1(n1187), .B0(a_s1[8]), .C0(n948), 
        .Y(n949) );
  OAI222_X0P5M_A12TR U1260 ( .A0(n949), .A1(n1358), .B0(n949), .B1(b_s1[19]), 
        .C0(n1189), .C1(n1204), .Y(n950) );
  AOI211_X0P5M_A12TR U1261 ( .A0(n1194), .A1(n1209), .B0(n951), .C0(n950), .Y(
        n999) );
  ADDF_X1M_A12TR U1262 ( .A(n954), .B(n953), .CI(n952), .CO(n1007), .S(n945)
         );
  OAI22_X0P5M_A12TR U1263 ( .A0(n1217), .A1(n1200), .B0(n1221), .B1(n1198), 
        .Y(n958) );
  AOI22_X0P5M_A12TR U1264 ( .A0(b_s1[18]), .A1(n1328), .B0(n1325), .B1(n1214), 
        .Y(n955) );
  OAI211_X0P5M_A12TR U1265 ( .A0(n1203), .A1(n1217), .B0(a_s1[11]), .C0(n955), 
        .Y(n956) );
  AOI211_X0P5M_A12TR U1266 ( .A0(n1210), .A1(n1214), .B0(n958), .C0(n957), .Y(
        n1006) );
  ADDF_X1M_A12TR U1267 ( .A(n961), .B(n960), .CI(n959), .CO(n1014), .S(n952)
         );
  INV_X0P5B_A12TR U1268 ( .A(n1233), .Y(n1230) );
  OAI22_X0P5M_A12TR U1269 ( .A0(n1235), .A1(n1216), .B0(n1215), .B1(n1230), 
        .Y(n965) );
  AOI22_X0P5M_A12TR U1270 ( .A0(n1304), .A1(b_s1[13]), .B0(n1308), .B1(
        b_s1[14]), .Y(n962) );
  OAI211_X0P5M_A12TR U1271 ( .A0(n1230), .A1(n1219), .B0(a_s1[14]), .C0(n962), 
        .Y(n963) );
  OAI222_X0P5M_A12TR U1272 ( .A0(n963), .A1(n1307), .B0(n963), .B1(b_s1[15]), 
        .C0(n1222), .C1(n1237), .Y(n964) );
  AOI211_X0P5M_A12TR U1273 ( .A0(b_s1[13]), .A1(n1226), .B0(n965), .C0(n964), 
        .Y(n1013) );
  ADDF_X1M_A12TR U1274 ( .A(n968), .B(n967), .CI(n966), .CO(n1022), .S(n959)
         );
  OAI22_X0P5M_A12TR U1275 ( .A0(n971), .A1(n1232), .B0(n1231), .B1(n969), .Y(
        n974) );
  AOI22_X0P5M_A12TR U1276 ( .A0(b_s1[10]), .A1(n1336), .B0(n1334), .B1(n1267), 
        .Y(n970) );
  OAI211_X0P5M_A12TR U1277 ( .A0(n1236), .A1(n971), .B0(a_s1[17]), .C0(n970), 
        .Y(n972) );
  AOI211_X0P5M_A12TR U1278 ( .A0(b_s1[10]), .A1(n1242), .B0(n974), .C0(n973), 
        .Y(n1021) );
  INV_X0P5B_A12TR U1279 ( .A(a_s1[26]), .Y(n1420) );
  INV_X0P5B_A12TR U1280 ( .A(n1107), .Y(n1029) );
  NAND2_X0P5A_A12TR U1281 ( .A(b_s1[0]), .B(n1029), .Y(n1102) );
  AOI22_X0P5M_A12TR U1282 ( .A0(n1243), .A1(n1377), .B0(b_s1[1]), .B1(n1379), 
        .Y(n977) );
  AOI22_X0P5M_A12TR U1283 ( .A0(b_s1[3]), .A1(n1380), .B0(b_s1[2]), .B1(n1381), 
        .Y(n976) );
  NAND3_X0P5M_A12TR U1284 ( .A(n976), .B(n977), .C(a_s1[26]), .Y(n975) );
  AO21A1AI2_X0P5M_A12TR U1285 ( .A0(n977), .A1(n976), .B0(a_s1[26]), .C0(n975), 
        .Y(n1031) );
  XNOR3_X0P5M_A12TR U1286 ( .A(n1102), .B(n1032), .C(n1031), .Y(n1038) );
  ADDF_X1M_A12TR U1287 ( .A(n980), .B(n979), .CI(n978), .CO(n1037), .S(n986)
         );
  AOI22_X0P5M_A12TR U1288 ( .A0(b_s1[4]), .A1(n1330), .B0(b_s1[6]), .B1(n1329), 
        .Y(n983) );
  AOI22_X0P5M_A12TR U1289 ( .A0(b_s1[5]), .A1(n1333), .B0(n1331), .B1(n1253), 
        .Y(n982) );
  NAND3_X0P5M_A12TR U1290 ( .A(n982), .B(n983), .C(n1424), .Y(n981) );
  AO21A1AI2_X0P5M_A12TR U1291 ( .A0(n983), .A1(n982), .B0(n1424), .C0(n981), 
        .Y(n1036) );
  ADDF_X1M_A12TR U1292 ( .A(n986), .B(n985), .CI(n984), .CO(n1043), .S(n966)
         );
  AOI22_X0P5M_A12TR U1293 ( .A0(b_s1[7]), .A1(n1313), .B0(n1311), .B1(n1260), 
        .Y(n989) );
  AOI22_X0P5M_A12TR U1294 ( .A0(n1310), .A1(b_s1[8]), .B0(n1309), .B1(b_s1[9]), 
        .Y(n988) );
  NAND3_X0P5M_A12TR U1295 ( .A(n988), .B(n989), .C(n1383), .Y(n987) );
  AO21A1AI2_X0P5M_A12TR U1296 ( .A0(n989), .A1(n988), .B0(n1383), .C0(n987), 
        .Y(n1042) );
  NOR2_X0P5B_A12TR U1297 ( .A(reset), .B(n990), .Y(\outreg_stage2/N30 ) );
  ADDF_X1M_A12TR U1298 ( .A(n993), .B(n992), .CI(n991), .CO(n1060), .S(n1053)
         );
  OAI22_X0P5M_A12TR U1299 ( .A0(n1168), .A1(n1183), .B0(n1167), .B1(n1172), 
        .Y(n997) );
  AOI22_X0P5M_A12TR U1300 ( .A0(n1301), .A1(n1360), .B0(n1302), .B1(b_s1[25]), 
        .Y(n994) );
  OAI211_X0P5M_A12TR U1301 ( .A0(n1183), .A1(n1170), .B0(a_s1[5]), .C0(n994), 
        .Y(n995) );
  OAI222_X0P5M_A12TR U1302 ( .A0(n995), .A1(n1299), .B0(n995), .B1(b_s1[23]), 
        .C0(n1173), .C1(n1186), .Y(n996) );
  AOI211_X0P5M_A12TR U1303 ( .A0(n1178), .A1(n1360), .B0(n997), .C0(n996), .Y(
        n1059) );
  ADDF_X1M_A12TR U1304 ( .A(n1000), .B(n999), .CI(n998), .CO(n1068), .S(n991)
         );
  OAI22_X0P5M_A12TR U1305 ( .A0(n1188), .A1(n1182), .B0(n1199), .B1(n1184), 
        .Y(n1004) );
  AOI22_X0P5M_A12TR U1306 ( .A0(n1359), .A1(n1326), .B0(n1362), .B1(b_s1[22]), 
        .Y(n1001) );
  OAI211_X0P5M_A12TR U1307 ( .A0(n1199), .A1(n1187), .B0(a_s1[8]), .C0(n1001), 
        .Y(n1002) );
  OAI222_X0P5M_A12TR U1308 ( .A0(n1002), .A1(n1358), .B0(n1002), .B1(b_s1[20]), 
        .C0(n1189), .C1(n1202), .Y(n1003) );
  AOI211_X0P5M_A12TR U1309 ( .A0(n1326), .A1(n1194), .B0(n1004), .C0(n1003), 
        .Y(n1067) );
  ADDF_X1M_A12TR U1310 ( .A(n1007), .B(n1006), .CI(n1005), .CO(n1076), .S(n998) );
  OAI22_X0P5M_A12TR U1311 ( .A0(n1221), .A1(n1200), .B0(n1204), .B1(n1198), 
        .Y(n1011) );
  AOI22_X0P5M_A12TR U1312 ( .A0(n1306), .A1(n1325), .B0(b_s1[19]), .B1(n1328), 
        .Y(n1008) );
  OAI211_X0P5M_A12TR U1313 ( .A0(n1203), .A1(n1221), .B0(a_s1[11]), .C0(n1008), 
        .Y(n1009) );
  AOI211_X0P5M_A12TR U1314 ( .A0(n1306), .A1(n1210), .B0(n1011), .C0(n1010), 
        .Y(n1075) );
  ADDF_X1M_A12TR U1315 ( .A(n1014), .B(n1013), .CI(n1012), .CO(n1084), .S(
        n1005) );
  INV_X0P5B_A12TR U1316 ( .A(n1335), .Y(n1016) );
  OAI22_X0P5M_A12TR U1317 ( .A0(n1016), .A1(n1215), .B0(n1237), .B1(n1216), 
        .Y(n1019) );
  AOI22_X0P5M_A12TR U1318 ( .A0(n1304), .A1(b_s1[14]), .B0(n1308), .B1(
        b_s1[15]), .Y(n1015) );
  OAI211_X0P5M_A12TR U1319 ( .A0(n1016), .A1(n1219), .B0(a_s1[14]), .C0(n1015), 
        .Y(n1017) );
  OAI222_X0P5M_A12TR U1320 ( .A0(n1017), .A1(n1307), .B0(n1017), .B1(b_s1[16]), 
        .C0(n1222), .C1(n1086), .Y(n1018) );
  AOI211_X0P5M_A12TR U1321 ( .A0(b_s1[14]), .A1(n1226), .B0(n1019), .C0(n1018), 
        .Y(n1083) );
  ADDF_X1M_A12TR U1322 ( .A(n1022), .B(n1021), .CI(n1020), .CO(n1094), .S(
        n1012) );
  OAI22_X0P5M_A12TR U1323 ( .A0(n1023), .A1(n1231), .B0(n1025), .B1(n1232), 
        .Y(n1028) );
  AOI22_X0P5M_A12TR U1324 ( .A0(b_s1[11]), .A1(n1336), .B0(n1312), .B1(n1334), 
        .Y(n1024) );
  OAI211_X0P5M_A12TR U1325 ( .A0(n1236), .A1(n1025), .B0(a_s1[17]), .C0(n1024), 
        .Y(n1026) );
  AOI211_X0P5M_A12TR U1326 ( .A0(b_s1[11]), .A1(n1242), .B0(n1028), .C0(n1027), 
        .Y(n1093) );
  AND2_X0P5M_A12TR U1327 ( .A(n1106), .B(n1029), .Y(n1339) );
  XNOR2_X0P5M_A12TR U1328 ( .A(a_s1[28]), .B(a_s1[27]), .Y(n1108) );
  NOR2_X0P5B_A12TR U1329 ( .A(n1029), .B(n1108), .Y(n1340) );
  NOR2_X0P5B_A12TR U1330 ( .A(n1106), .B(n1107), .Y(n1341) );
  AOI222_X0P5M_A12TR U1331 ( .A0(b_s1[1]), .A1(n1339), .B0(b_s1[0]), .B1(n1340), .C0(n1298), .C1(n1341), .Y(n1103) );
  INV_X0P5B_A12TR U1332 ( .A(a_s1[29]), .Y(n1419) );
  OAI21_X0P5M_A12TR U1333 ( .A0(n1102), .A1(n1419), .B0(n1103), .Y(n1030) );
  OAI31_X0P5M_A12TR U1334 ( .A0(n1102), .A1(n1103), .A2(n1419), .B0(n1030), 
        .Y(n1117) );
  AO21B_X0P5M_A12TR U1335 ( .A0(n1102), .A1(n1032), .B0N(n1031), .Y(n1116) );
  AOI22_X0P5M_A12TR U1336 ( .A0(b_s1[2]), .A1(n1379), .B0(n1342), .B1(n1377), 
        .Y(n1035) );
  AOI22_X0P5M_A12TR U1337 ( .A0(b_s1[3]), .A1(n1381), .B0(b_s1[4]), .B1(n1380), 
        .Y(n1034) );
  NAND3_X0P5M_A12TR U1338 ( .A(n1034), .B(n1035), .C(n1420), .Y(n1033) );
  AO21A1AI2_X0P5M_A12TR U1339 ( .A0(n1035), .A1(n1034), .B0(n1420), .C0(n1033), 
        .Y(n1115) );
  ADDF_X1M_A12TR U1340 ( .A(n1038), .B(n1037), .CI(n1036), .CO(n1123), .S(
        n1044) );
  AOI22_X0P5M_A12TR U1341 ( .A0(b_s1[5]), .A1(n1330), .B0(b_s1[7]), .B1(n1329), 
        .Y(n1041) );
  AOI22_X0P5M_A12TR U1342 ( .A0(n1378), .A1(n1331), .B0(b_s1[6]), .B1(n1333), 
        .Y(n1040) );
  NAND3_X0P5M_A12TR U1343 ( .A(n1040), .B(n1041), .C(n1424), .Y(n1039) );
  AO21A1AI2_X0P5M_A12TR U1344 ( .A0(n1041), .A1(n1040), .B0(n1424), .C0(n1039), 
        .Y(n1122) );
  ADDF_X1M_A12TR U1345 ( .A(n1044), .B(n1043), .CI(n1042), .CO(n1130), .S(
        n1020) );
  AOI22_X0P5M_A12TR U1346 ( .A0(n1313), .A1(b_s1[8]), .B0(n1311), .B1(n1332), 
        .Y(n1047) );
  AOI22_X0P5M_A12TR U1347 ( .A0(n1310), .A1(b_s1[9]), .B0(n1309), .B1(b_s1[10]), .Y(n1046) );
  NAND3_X0P5M_A12TR U1348 ( .A(n1046), .B(n1047), .C(n1383), .Y(n1045) );
  AO21A1AI2_X0P5M_A12TR U1349 ( .A0(n1047), .A1(n1046), .B0(n1383), .C0(n1045), 
        .Y(n1129) );
  ADDF_X1M_A12TR U1350 ( .A(b_s1[26]), .B(b_s1[27]), .CI(n1048), .CO(n1136), 
        .S(n1177) );
  INV_X0P5B_A12TR U1351 ( .A(b_s1[27]), .Y(n1166) );
  AOI22_X0P5M_A12TR U1352 ( .A0(n1376), .A1(b_s1[26]), .B0(b_s1[28]), .B1(
        n1375), .Y(n1049) );
  OAI211_X0P5M_A12TR U1353 ( .A0(n1166), .A1(n1370), .B0(a_s1[2]), .C0(n1049), 
        .Y(n1051) );
  AOI22_X0P5M_A12TR U1354 ( .A0(n1157), .A1(n1300), .B0(n1156), .B1(b_s1[28]), 
        .Y(n1050) );
  AO21A1AI2_X0P5M_A12TR U1355 ( .A0(n1300), .A1(n1373), .B0(n1051), .C0(n1050), 
        .Y(n1052) );
  AOI21_X0P5M_A12TR U1356 ( .A0(n1162), .A1(b_s1[27]), .B0(n1052), .Y(n1145)
         );
  ADDF_X1M_A12TR U1357 ( .A(n1055), .B(n1054), .CI(n1053), .CO(n1144), .S(n990) );
  XNOR2_X0P5M_A12TR U1358 ( .A(n1145), .B(n1144), .Y(n1057) );
  OAI21_X0P5M_A12TR U1359 ( .A0(n1146), .A1(n1057), .B0(n1450), .Y(n1056) );
  AOI21_X0P5M_A12TR U1360 ( .A0(n1146), .A1(n1057), .B0(n1056), .Y(
        \outreg_stage2/N31 ) );
  ADDF_X1M_A12TR U1361 ( .A(n1060), .B(n1059), .CI(n1058), .CO(n1165), .S(
        n1146) );
  OAI22_X0P5M_A12TR U1362 ( .A0(n1168), .A1(n1172), .B0(n1167), .B1(n1171), 
        .Y(n1064) );
  AOI22_X0P5M_A12TR U1363 ( .A0(n1301), .A1(n1065), .B0(n1302), .B1(b_s1[26]), 
        .Y(n1061) );
  OAI211_X0P5M_A12TR U1364 ( .A0(n1172), .A1(n1170), .B0(a_s1[5]), .C0(n1061), 
        .Y(n1062) );
  OAI222_X0P5M_A12TR U1365 ( .A0(n1062), .A1(n1299), .B0(n1062), .B1(b_s1[24]), 
        .C0(n1173), .C1(n1183), .Y(n1063) );
  AOI211_X0P5M_A12TR U1366 ( .A0(n1178), .A1(n1065), .B0(n1064), .C0(n1063), 
        .Y(n1164) );
  ADDF_X1M_A12TR U1367 ( .A(n1068), .B(n1067), .CI(n1066), .CO(n1181), .S(
        n1058) );
  OAI22_X0P5M_A12TR U1368 ( .A0(n1186), .A1(n1182), .B0(n1188), .B1(n1184), 
        .Y(n1072) );
  AOI22_X0P5M_A12TR U1369 ( .A0(n1359), .A1(n1073), .B0(b_s1[23]), .B1(n1362), 
        .Y(n1069) );
  OAI211_X0P5M_A12TR U1370 ( .A0(n1188), .A1(n1187), .B0(a_s1[8]), .C0(n1069), 
        .Y(n1070) );
  OAI222_X0P5M_A12TR U1371 ( .A0(n1070), .A1(n1358), .B0(n1070), .B1(b_s1[21]), 
        .C0(n1189), .C1(n1199), .Y(n1071) );
  AOI211_X0P5M_A12TR U1372 ( .A0(n1194), .A1(n1073), .B0(n1072), .C0(n1071), 
        .Y(n1180) );
  ADDF_X1M_A12TR U1373 ( .A(n1076), .B(n1075), .CI(n1074), .CO(n1197), .S(
        n1066) );
  OAI22_X0P5M_A12TR U1374 ( .A0(n1204), .A1(n1200), .B0(n1202), .B1(n1198), 
        .Y(n1080) );
  AOI22_X0P5M_A12TR U1375 ( .A0(n1325), .A1(n1081), .B0(b_s1[20]), .B1(n1328), 
        .Y(n1077) );
  OAI211_X0P5M_A12TR U1376 ( .A0(n1203), .A1(n1204), .B0(a_s1[11]), .C0(n1077), 
        .Y(n1078) );
  AOI211_X0P5M_A12TR U1377 ( .A0(n1210), .A1(n1081), .B0(n1080), .C0(n1079), 
        .Y(n1196) );
  ADDF_X1M_A12TR U1378 ( .A(n1084), .B(n1083), .CI(n1082), .CO(n1213), .S(
        n1074) );
  INV_X0P5B_A12TR U1379 ( .A(n1085), .Y(n1088) );
  OAI22_X0P5M_A12TR U1380 ( .A0(n1086), .A1(n1216), .B0(n1215), .B1(n1088), 
        .Y(n1091) );
  AOI22_X0P5M_A12TR U1381 ( .A0(n1304), .A1(b_s1[15]), .B0(n1308), .B1(
        b_s1[16]), .Y(n1087) );
  OAI211_X0P5M_A12TR U1382 ( .A0(n1088), .A1(n1219), .B0(a_s1[14]), .C0(n1087), 
        .Y(n1089) );
  OAI222_X0P5M_A12TR U1383 ( .A0(n1089), .A1(n1307), .B0(n1089), .B1(b_s1[17]), 
        .C0(n1222), .C1(n1217), .Y(n1090) );
  AOI211_X0P5M_A12TR U1384 ( .A0(b_s1[15]), .A1(n1226), .B0(n1091), .C0(n1090), 
        .Y(n1212) );
  ADDF_X1M_A12TR U1385 ( .A(n1094), .B(n1093), .CI(n1092), .CO(n1229), .S(
        n1082) );
  OAI22_X0P5M_A12TR U1386 ( .A0(n1098), .A1(n1232), .B0(n1231), .B1(n1095), 
        .Y(n1101) );
  AOI22_X0P5M_A12TR U1387 ( .A0(b_s1[12]), .A1(n1336), .B0(n1334), .B1(n1096), 
        .Y(n1097) );
  OAI211_X0P5M_A12TR U1388 ( .A0(n1236), .A1(n1098), .B0(a_s1[17]), .C0(n1097), 
        .Y(n1099) );
  AOI211_X0P5M_A12TR U1389 ( .A0(b_s1[12]), .A1(n1242), .B0(n1101), .C0(n1100), 
        .Y(n1228) );
  INV_X0P5B_A12TR U1390 ( .A(n1102), .Y(n1105) );
  NAND2_X0P5A_A12TR U1391 ( .A(a_s1[29]), .B(n1103), .Y(n1104) );
  NOR2_X0P5B_A12TR U1392 ( .A(n1105), .B(n1104), .Y(n1114) );
  NOR3BB_X0P5M_A12TR U1393 ( .AN(n1108), .BN(n1107), .C(n1106), .Y(n1343) );
  AOI22_X0P5M_A12TR U1394 ( .A0(b_s1[0]), .A1(n1343), .B0(n1109), .B1(n1341), 
        .Y(n1112) );
  AOI22_X0P5M_A12TR U1395 ( .A0(b_s1[1]), .A1(n1340), .B0(b_s1[2]), .B1(n1339), 
        .Y(n1111) );
  NAND3_X0P5M_A12TR U1396 ( .A(n1111), .B(n1112), .C(a_s1[29]), .Y(n1110) );
  AO21A1AI2_X0P5M_A12TR U1397 ( .A0(n1112), .A1(n1111), .B0(a_s1[29]), .C0(
        n1110), .Y(n1113) );
  NAND2_X0P5A_A12TR U1398 ( .A(n1114), .B(n1113), .Y(n1248) );
  OAI21_X0P5M_A12TR U1399 ( .A0(n1114), .A1(n1113), .B0(n1248), .Y(n1252) );
  ADDF_X1M_A12TR U1400 ( .A(n1117), .B(n1116), .CI(n1115), .CO(n1251), .S(
        n1124) );
  AOI22_X0P5M_A12TR U1401 ( .A0(b_s1[3]), .A1(n1379), .B0(n1118), .B1(n1377), 
        .Y(n1121) );
  AOI22_X0P5M_A12TR U1402 ( .A0(b_s1[4]), .A1(n1381), .B0(b_s1[5]), .B1(n1380), 
        .Y(n1120) );
  NAND3_X0P5M_A12TR U1403 ( .A(n1120), .B(n1121), .C(n1420), .Y(n1119) );
  AO21A1AI2_X0P5M_A12TR U1404 ( .A0(n1121), .A1(n1120), .B0(n1420), .C0(n1119), 
        .Y(n1250) );
  ADDF_X1M_A12TR U1405 ( .A(n1124), .B(n1123), .CI(n1122), .CO(n1258), .S(
        n1131) );
  AOI22_X0P5M_A12TR U1406 ( .A0(b_s1[6]), .A1(n1330), .B0(b_s1[8]), .B1(n1329), 
        .Y(n1128) );
  AOI22_X0P5M_A12TR U1407 ( .A0(b_s1[7]), .A1(n1333), .B0(n1331), .B1(n1125), 
        .Y(n1127) );
  NAND3_X0P5M_A12TR U1408 ( .A(n1127), .B(n1128), .C(n1424), .Y(n1126) );
  AO21A1AI2_X0P5M_A12TR U1409 ( .A0(n1128), .A1(n1127), .B0(n1424), .C0(n1126), 
        .Y(n1257) );
  ADDF_X1M_A12TR U1410 ( .A(n1131), .B(n1130), .CI(n1129), .CO(n1265), .S(
        n1092) );
  AOI22_X0P5M_A12TR U1411 ( .A0(n1313), .A1(b_s1[9]), .B0(n1311), .B1(n1132), 
        .Y(n1135) );
  AOI22_X0P5M_A12TR U1412 ( .A0(b_s1[11]), .A1(n1309), .B0(n1310), .B1(
        b_s1[10]), .Y(n1134) );
  NAND3_X0P5M_A12TR U1413 ( .A(n1134), .B(n1135), .C(n1383), .Y(n1133) );
  AO21A1AI2_X0P5M_A12TR U1414 ( .A0(n1135), .A1(n1134), .B0(n1383), .C0(n1133), 
        .Y(n1264) );
  ADDF_X1M_A12TR U1415 ( .A(b_s1[27]), .B(b_s1[28]), .CI(n1136), .CO(n1153), 
        .S(n1300) );
  INV_X0P5B_A12TR U1416 ( .A(b_s1[28]), .Y(n1138) );
  AOI22_X0P5M_A12TR U1417 ( .A0(n1376), .A1(b_s1[27]), .B0(b_s1[29]), .B1(
        n1375), .Y(n1137) );
  OAI211_X0P5M_A12TR U1418 ( .A0(n1138), .A1(n1370), .B0(a_s1[2]), .C0(n1137), 
        .Y(n1140) );
  AOI22_X0P5M_A12TR U1419 ( .A0(n1157), .A1(n1142), .B0(n1156), .B1(b_s1[29]), 
        .Y(n1139) );
  AO21A1AI2_X0P5M_A12TR U1420 ( .A0(n1142), .A1(n1141), .B0(n1140), .C0(n1139), 
        .Y(n1143) );
  AOI21_X0P5M_A12TR U1421 ( .A0(n1162), .A1(b_s1[28]), .B0(n1143), .Y(n1150)
         );
  XOR2_X0P5M_A12TR U1422 ( .A(n1151), .B(n1150), .Y(n1148) );
  CGENI_X1M_A12TR U1423 ( .A(n1146), .B(n1145), .CI(n1144), .CON(n1149) );
  OAI21_X0P5M_A12TR U1424 ( .A0(n1148), .A1(n1149), .B0(n1450), .Y(n1147) );
  AOI21_X0P5M_A12TR U1425 ( .A0(n1148), .A1(n1149), .B0(n1147), .Y(
        \outreg_stage2/N32 ) );
  INV_X0P5B_A12TR U1426 ( .A(n1149), .Y(n1152) );
  CGEN_X1M_A12TR U1427 ( .A(n1152), .B(n1151), .CI(n1150), .CO(n1397) );
  ADDF_X1M_A12TR U1428 ( .A(b_s1[28]), .B(b_s1[29]), .CI(n1153), .CO(n1368), 
        .S(n1142) );
  INV_X0P5B_A12TR U1429 ( .A(b_s1[29]), .Y(n1155) );
  AOI22_X0P5M_A12TR U1430 ( .A0(n1376), .A1(b_s1[28]), .B0(b_s1[30]), .B1(
        n1375), .Y(n1154) );
  OAI211_X0P5M_A12TR U1431 ( .A0(n1155), .A1(n1370), .B0(a_s1[2]), .C0(n1154), 
        .Y(n1159) );
  AOI22_X0P5M_A12TR U1432 ( .A0(n1157), .A1(n1160), .B0(n1156), .B1(b_s1[30]), 
        .Y(n1158) );
  AO21A1AI2_X0P5M_A12TR U1433 ( .A0(n1160), .A1(n1373), .B0(n1159), .C0(n1158), 
        .Y(n1161) );
  AOI21_X0P5M_A12TR U1434 ( .A0(n1162), .A1(b_s1[29]), .B0(n1161), .Y(n1396)
         );
  ADDF_X1M_A12TR U1435 ( .A(n1165), .B(n1164), .CI(n1163), .CO(n1394), .S(
        n1151) );
  OAI22_X0P5M_A12TR U1436 ( .A0(n1168), .A1(n1171), .B0(n1167), .B1(n1166), 
        .Y(n1176) );
  AOI22_X0P5M_A12TR U1437 ( .A0(n1301), .A1(n1177), .B0(n1302), .B1(b_s1[27]), 
        .Y(n1169) );
  OAI211_X0P5M_A12TR U1438 ( .A0(n1171), .A1(n1170), .B0(a_s1[5]), .C0(n1169), 
        .Y(n1174) );
  OAI222_X0P5M_A12TR U1439 ( .A0(n1174), .A1(n1299), .B0(n1174), .B1(b_s1[25]), 
        .C0(n1173), .C1(n1172), .Y(n1175) );
  AOI211_X0P5M_A12TR U1440 ( .A0(n1178), .A1(n1177), .B0(n1176), .C0(n1175), 
        .Y(n1393) );
  ADDF_X1M_A12TR U1441 ( .A(n1181), .B(n1180), .CI(n1179), .CO(n1409), .S(
        n1163) );
  OAI22_X0P5M_A12TR U1442 ( .A0(n1186), .A1(n1184), .B0(n1183), .B1(n1182), 
        .Y(n1192) );
  AOI22_X0P5M_A12TR U1443 ( .A0(n1359), .A1(n1193), .B0(n1362), .B1(b_s1[24]), 
        .Y(n1185) );
  OAI211_X0P5M_A12TR U1444 ( .A0(n1187), .A1(n1186), .B0(a_s1[8]), .C0(n1185), 
        .Y(n1190) );
  OAI222_X0P5M_A12TR U1445 ( .A0(n1190), .A1(n1358), .B0(n1190), .B1(b_s1[22]), 
        .C0(n1189), .C1(n1188), .Y(n1191) );
  AOI211_X0P5M_A12TR U1446 ( .A0(n1194), .A1(n1193), .B0(n1192), .C0(n1191), 
        .Y(n1408) );
  ADDF_X1M_A12TR U1447 ( .A(n1197), .B(n1196), .CI(n1195), .CO(n1391), .S(
        n1179) );
  OAI22_X0P5M_A12TR U1448 ( .A0(n1202), .A1(n1200), .B0(n1199), .B1(n1198), 
        .Y(n1208) );
  AOI22_X0P5M_A12TR U1449 ( .A0(n1325), .A1(n1209), .B0(n1328), .B1(b_s1[21]), 
        .Y(n1201) );
  OAI211_X0P5M_A12TR U1450 ( .A0(n1203), .A1(n1202), .B0(a_s1[11]), .C0(n1201), 
        .Y(n1206) );
  OAI222_X0P5M_A12TR U1451 ( .A0(n1206), .A1(n1324), .B0(n1206), .B1(b_s1[19]), 
        .C0(n1205), .C1(n1204), .Y(n1207) );
  AOI211_X0P5M_A12TR U1452 ( .A0(n1210), .A1(n1209), .B0(n1208), .C0(n1207), 
        .Y(n1390) );
  ADDF_X1M_A12TR U1453 ( .A(n1213), .B(n1212), .CI(n1211), .CO(n1418), .S(
        n1195) );
  INV_X0P5B_A12TR U1454 ( .A(n1214), .Y(n1220) );
  OAI22_X0P5M_A12TR U1455 ( .A0(n1217), .A1(n1216), .B0(n1215), .B1(n1220), 
        .Y(n1225) );
  AOI22_X0P5M_A12TR U1456 ( .A0(n1304), .A1(b_s1[16]), .B0(b_s1[17]), .B1(
        n1308), .Y(n1218) );
  OAI211_X0P5M_A12TR U1457 ( .A0(n1220), .A1(n1219), .B0(a_s1[14]), .C0(n1218), 
        .Y(n1223) );
  OAI222_X0P5M_A12TR U1458 ( .A0(n1223), .A1(n1307), .B0(n1223), .B1(b_s1[18]), 
        .C0(n1222), .C1(n1221), .Y(n1224) );
  AOI211_X0P5M_A12TR U1459 ( .A0(b_s1[16]), .A1(n1226), .B0(n1225), .C0(n1224), 
        .Y(n1417) );
  ADDF_X1M_A12TR U1460 ( .A(n1229), .B(n1228), .CI(n1227), .CO(n1412), .S(
        n1211) );
  OAI22_X0P5M_A12TR U1461 ( .A0(n1235), .A1(n1232), .B0(n1231), .B1(n1230), 
        .Y(n1241) );
  AOI22_X0P5M_A12TR U1462 ( .A0(b_s1[13]), .A1(n1336), .B0(n1334), .B1(n1233), 
        .Y(n1234) );
  OAI211_X0P5M_A12TR U1463 ( .A0(n1236), .A1(n1235), .B0(a_s1[17]), .C0(n1234), 
        .Y(n1239) );
  AOI211_X0P5M_A12TR U1464 ( .A0(b_s1[13]), .A1(n1242), .B0(n1241), .C0(n1240), 
        .Y(n1411) );
  AOI22_X0P5M_A12TR U1465 ( .A0(n1243), .A1(n1341), .B0(b_s1[1]), .B1(n1343), 
        .Y(n1246) );
  AOI22_X0P5M_A12TR U1466 ( .A0(b_s1[3]), .A1(n1339), .B0(b_s1[2]), .B1(n1340), 
        .Y(n1245) );
  NAND3_X0P5M_A12TR U1467 ( .A(n1245), .B(n1246), .C(a_s1[29]), .Y(n1244) );
  AO21A1AI2_X0P5M_A12TR U1468 ( .A0(n1246), .A1(n1245), .B0(a_s1[29]), .C0(
        n1244), .Y(n1452) );
  INV_X0P5B_A12TR U1469 ( .A(n1297), .Y(n1293) );
  OAI21_X0P5M_A12TR U1470 ( .A0(n1247), .A1(n1293), .B0(n1248), .Y(n1453) );
  OAI31_X0P5M_A12TR U1471 ( .A0(n1248), .A1(n1247), .A2(n1293), .B0(n1453), 
        .Y(n1249) );
  XOR2_X0P5M_A12TR U1472 ( .A(n1452), .B(n1249), .Y(n1403) );
  ADDF_X1M_A12TR U1473 ( .A(n1252), .B(n1251), .CI(n1250), .CO(n1402), .S(
        n1259) );
  AOI22_X0P5M_A12TR U1474 ( .A0(b_s1[4]), .A1(n1379), .B0(n1377), .B1(n1253), 
        .Y(n1256) );
  AOI22_X0P5M_A12TR U1475 ( .A0(b_s1[5]), .A1(n1381), .B0(b_s1[6]), .B1(n1380), 
        .Y(n1255) );
  NAND3_X0P5M_A12TR U1476 ( .A(n1255), .B(n1256), .C(n1420), .Y(n1254) );
  AO21A1AI2_X0P5M_A12TR U1477 ( .A0(n1256), .A1(n1255), .B0(n1420), .C0(n1254), 
        .Y(n1401) );
  ADDF_X1M_A12TR U1478 ( .A(n1259), .B(n1258), .CI(n1257), .CO(n1387), .S(
        n1266) );
  AOI22_X0P5M_A12TR U1479 ( .A0(b_s1[7]), .A1(n1330), .B0(n1329), .B1(b_s1[9]), 
        .Y(n1263) );
  AOI22_X0P5M_A12TR U1480 ( .A0(b_s1[8]), .A1(n1333), .B0(n1331), .B1(n1260), 
        .Y(n1262) );
  NAND3_X0P5M_A12TR U1481 ( .A(n1262), .B(n1263), .C(n1424), .Y(n1261) );
  AO21A1AI2_X0P5M_A12TR U1482 ( .A0(n1263), .A1(n1262), .B0(n1424), .C0(n1261), 
        .Y(n1386) );
  ADDF_X1M_A12TR U1483 ( .A(n1266), .B(n1265), .CI(n1264), .CO(n1405), .S(
        n1227) );
  AOI22_X0P5M_A12TR U1484 ( .A0(n1313), .A1(b_s1[10]), .B0(n1311), .B1(n1267), 
        .Y(n1270) );
  AOI22_X0P5M_A12TR U1485 ( .A0(b_s1[11]), .A1(n1310), .B0(b_s1[12]), .B1(
        n1309), .Y(n1269) );
  NAND3_X0P5M_A12TR U1486 ( .A(n1269), .B(n1270), .C(n1383), .Y(n1268) );
  AO21A1AI2_X0P5M_A12TR U1487 ( .A0(n1270), .A1(n1269), .B0(n1383), .C0(n1268), 
        .Y(n1404) );
  NOR2_X0P5B_A12TR U1488 ( .A(reset), .B(n1271), .Y(\outreg_stage2/N33 ) );
  NAND2_X0P5A_A12TR U1489 ( .A(a_s1[0]), .B(b_s1[0]), .Y(n1275) );
  NOR2_X0P5B_A12TR U1490 ( .A(reset), .B(n1275), .Y(\outreg_stage2/N3 ) );
  OAI31_X0P5M_A12TR U1491 ( .A0(n1425), .A1(n1274), .A2(n1275), .B0(n1450), 
        .Y(n1273) );
  OA21A1OI2_X0P7M_A12TR U1492 ( .A0(n1425), .A1(n1275), .B0(n1274), .C0(n1273), 
        .Y(\outreg_stage2/N4 ) );
  OA211_X0P5M_A12TR U1493 ( .A0(n1277), .A1(n1276), .B0(n1450), .C0(n1278), 
        .Y(\outreg_stage2/N5 ) );
  XOR2_X0P5M_A12TR U1494 ( .A(n1279), .B(n1278), .Y(n1281) );
  NOR2_X0P5B_A12TR U1495 ( .A(n1282), .B(n1281), .Y(n1280) );
  XOR2_X0P5M_A12TR U1496 ( .A(n1284), .B(n1283), .Y(n1286) );
  NOR2_X0P5B_A12TR U1497 ( .A(n1287), .B(n1286), .Y(n1285) );
  XNOR2_X0P5M_A12TR U1498 ( .A(n1289), .B(n1288), .Y(n1291) );
  NOR2_X0P5B_A12TR U1499 ( .A(n1292), .B(n1291), .Y(n1290) );
  OAI211_X0P5M_A12TR U1500 ( .A0(a_s1[30]), .A1(a_s1[31]), .B0(b_s1[0]), .C0(
        n1293), .Y(n1295) );
  NAND2_X0P5A_A12TR U1501 ( .A(b_s1[1]), .B(n1297), .Y(n1294) );
  AOI31_X0P5M_A12TR U1502 ( .A0(n1298), .A1(n1297), .A2(a_s1[31]), .B0(n1296), 
        .Y(n1449) );
  AOI22_X0P5M_A12TR U1503 ( .A0(n1301), .A1(n1300), .B0(n1299), .B1(b_s1[26]), 
        .Y(n1323) );
  AOI22_X0P5M_A12TR U1504 ( .A0(n1303), .A1(b_s1[27]), .B0(n1302), .B1(
        b_s1[28]), .Y(n1322) );
  AOI22_X0P5M_A12TR U1505 ( .A0(n1306), .A1(n1305), .B0(n1304), .B1(b_s1[17]), 
        .Y(n1319) );
  AOI22_X0P5M_A12TR U1506 ( .A0(n1308), .A1(b_s1[18]), .B0(n1307), .B1(
        b_s1[19]), .Y(n1318) );
  AOI22_X0P5M_A12TR U1507 ( .A0(n1310), .A1(b_s1[12]), .B0(n1309), .B1(
        b_s1[13]), .Y(n1315) );
  AOI22_X0P5M_A12TR U1508 ( .A0(n1313), .A1(b_s1[11]), .B0(n1312), .B1(n1311), 
        .Y(n1314) );
  NAND2_X0P5A_A12TR U1509 ( .A(n1315), .B(n1314), .Y(n1317) );
  NAND3_X0P5M_A12TR U1510 ( .A(n1318), .B(n1319), .C(n1317), .Y(n1316) );
  AO21A1AI2_X0P5M_A12TR U1511 ( .A0(n1319), .A1(n1318), .B0(n1317), .C0(n1316), 
        .Y(n1321) );
  NAND3_X0P5M_A12TR U1512 ( .A(n1322), .B(n1323), .C(n1321), .Y(n1320) );
  AO21A1AI2_X0P5M_A12TR U1513 ( .A0(n1323), .A1(n1322), .B0(n1321), .C0(n1320), 
        .Y(n1367) );
  AOI22_X0P5M_A12TR U1514 ( .A0(n1326), .A1(n1325), .B0(n1324), .B1(b_s1[20]), 
        .Y(n1357) );
  AOI22_X0P5M_A12TR U1515 ( .A0(n1328), .A1(b_s1[22]), .B0(n1327), .B1(
        b_s1[21]), .Y(n1356) );
  AOI22_X0P5M_A12TR U1516 ( .A0(n1330), .A1(b_s1[8]), .B0(n1329), .B1(b_s1[10]), .Y(n1353) );
  AOI22_X0P5M_A12TR U1517 ( .A0(n1333), .A1(b_s1[9]), .B0(n1332), .B1(n1331), 
        .Y(n1352) );
  AOI22_X0P5M_A12TR U1518 ( .A0(n1336), .A1(b_s1[14]), .B0(n1335), .B1(n1334), 
        .Y(n1349) );
  AOI22_X0P5M_A12TR U1519 ( .A0(n1338), .A1(b_s1[15]), .B0(n1337), .B1(
        b_s1[16]), .Y(n1348) );
  AOI22_X0P5M_A12TR U1520 ( .A0(b_s1[3]), .A1(n1340), .B0(b_s1[4]), .B1(n1339), 
        .Y(n1345) );
  AOI22_X0P5M_A12TR U1521 ( .A0(b_s1[2]), .A1(n1343), .B0(n1342), .B1(n1341), 
        .Y(n1344) );
  NAND2_X0P5A_A12TR U1522 ( .A(n1345), .B(n1344), .Y(n1347) );
  NAND3_X0P5M_A12TR U1523 ( .A(n1348), .B(n1349), .C(n1347), .Y(n1346) );
  AO21A1AI2_X0P5M_A12TR U1524 ( .A0(n1349), .A1(n1348), .B0(n1347), .C0(n1346), 
        .Y(n1351) );
  NAND3_X0P5M_A12TR U1525 ( .A(n1352), .B(n1353), .C(n1351), .Y(n1350) );
  AO21A1AI2_X0P5M_A12TR U1526 ( .A0(n1353), .A1(n1352), .B0(n1351), .C0(n1350), 
        .Y(n1355) );
  NAND3_X0P5M_A12TR U1527 ( .A(n1356), .B(n1357), .C(n1355), .Y(n1354) );
  AO21A1AI2_X0P5M_A12TR U1528 ( .A0(n1357), .A1(n1356), .B0(n1355), .C0(n1354), 
        .Y(n1366) );
  AOI22_X0P5M_A12TR U1529 ( .A0(n1360), .A1(n1359), .B0(n1358), .B1(b_s1[23]), 
        .Y(n1364) );
  AOI22_X0P5M_A12TR U1530 ( .A0(n1362), .A1(b_s1[25]), .B0(n1361), .B1(
        b_s1[24]), .Y(n1363) );
  NAND2_X0P5A_A12TR U1531 ( .A(n1364), .B(n1363), .Y(n1365) );
  XOR3_X0P5M_A12TR U1532 ( .A(n1367), .B(n1366), .C(n1365), .Y(n1448) );
  ADDF_X1M_A12TR U1533 ( .A(b_s1[29]), .B(b_s1[30]), .CI(n1368), .CO(n1369), 
        .S(n1160) );
  XOR2_X0P5M_A12TR U1534 ( .A(b_s1[31]), .B(n1369), .Y(n1374) );
  AO21A1AI2_X0P5M_A12TR U1535 ( .A0(n1374), .A1(b_s1[30]), .B0(n1371), .C0(
        n1370), .Y(n1372) );
  AO21A1AI2_X0P5M_A12TR U1536 ( .A0(n1374), .A1(n1373), .B0(b_s1[30]), .C0(
        n1372), .Y(n1446) );
  AOI22_X0P5M_A12TR U1537 ( .A0(n1376), .A1(b_s1[29]), .B0(b_s1[31]), .B1(
        n1375), .Y(n1445) );
  AOI22_X0P5M_A12TR U1538 ( .A0(b_s1[5]), .A1(n1379), .B0(n1378), .B1(n1377), 
        .Y(n1442) );
  AOI22_X0P5M_A12TR U1539 ( .A0(n1381), .A1(b_s1[6]), .B0(n1380), .B1(b_s1[7]), 
        .Y(n1441) );
  AOI22_X0P5M_A12TR U1540 ( .A0(a_s1[17]), .A1(a_s1[20]), .B0(n1383), .B1(
        n1382), .Y(n1438) );
  AOI22_X0P5M_A12TR U1541 ( .A0(a_s1[8]), .A1(a_s1[14]), .B0(n1385), .B1(n1384), .Y(n1437) );
  ADDF_X1M_A12TR U1542 ( .A(n1388), .B(n1387), .CI(n1386), .CO(n1435), .S(
        n1406) );
  ADDF_X1M_A12TR U1543 ( .A(n1391), .B(n1390), .CI(n1389), .CO(n1400), .S(
        n1407) );
  ADDF_X1M_A12TR U1544 ( .A(n1394), .B(n1393), .CI(n1392), .CO(n1399), .S(
        n1395) );
  ADDF_X1M_A12TR U1545 ( .A(n1397), .B(n1396), .CI(n1395), .CO(n1398), .S(
        n1271) );
  XOR3_X0P5M_A12TR U1546 ( .A(n1400), .B(n1399), .C(n1398), .Y(n1434) );
  ADDF_X1M_A12TR U1547 ( .A(n1403), .B(n1402), .CI(n1401), .CO(n1432), .S(
        n1388) );
  ADDF_X1M_A12TR U1548 ( .A(n1406), .B(n1405), .CI(n1404), .CO(n1415), .S(
        n1410) );
  ADDF_X1M_A12TR U1549 ( .A(n1409), .B(n1408), .CI(n1407), .CO(n1414), .S(
        n1392) );
  ADDF_X1M_A12TR U1550 ( .A(n1412), .B(n1411), .CI(n1410), .CO(n1413), .S(
        n1416) );
  XOR3_X0P5M_A12TR U1551 ( .A(n1415), .B(n1414), .C(n1413), .Y(n1431) );
  ADDF_X1M_A12TR U1552 ( .A(n1418), .B(n1417), .CI(n1416), .CO(n1422), .S(
        n1389) );
  AOI22_X0P5M_A12TR U1553 ( .A0(a_s1[29]), .A1(a_s1[26]), .B0(n1420), .B1(
        n1419), .Y(n1421) );
  XNOR2_X0P5M_A12TR U1554 ( .A(n1422), .B(n1421), .Y(n1429) );
  AOI22_X0P5M_A12TR U1555 ( .A0(a_s1[5]), .A1(a_s1[23]), .B0(n1424), .B1(n1423), .Y(n1428) );
  AOI22_X0P5M_A12TR U1556 ( .A0(a_s1[2]), .A1(a_s1[11]), .B0(n1426), .B1(n1425), .Y(n1427) );
  XNOR3_X0P5M_A12TR U1557 ( .A(n1429), .B(n1428), .C(n1427), .Y(n1430) );
  XNOR3_X0P5M_A12TR U1558 ( .A(n1432), .B(n1431), .C(n1430), .Y(n1433) );
  XNOR3_X0P5M_A12TR U1559 ( .A(n1435), .B(n1434), .C(n1433), .Y(n1436) );
  XNOR3_X0P5M_A12TR U1560 ( .A(n1438), .B(n1437), .C(n1436), .Y(n1440) );
  NAND3_X0P5M_A12TR U1561 ( .A(n1441), .B(n1442), .C(n1440), .Y(n1439) );
  AO21A1AI2_X0P5M_A12TR U1562 ( .A0(n1442), .A1(n1441), .B0(n1440), .C0(n1439), 
        .Y(n1444) );
  NAND3_X0P5M_A12TR U1563 ( .A(n1445), .B(n1446), .C(n1444), .Y(n1443) );
  AO21A1AI2_X0P5M_A12TR U1564 ( .A0(n1446), .A1(n1445), .B0(n1444), .C0(n1443), 
        .Y(n1447) );
  XNOR3_X0P5M_A12TR U1565 ( .A(n1449), .B(n1448), .C(n1447), .Y(n1454) );
  AO21A1AI2_X0P5M_A12TR U1566 ( .A0(n1453), .A1(n1452), .B0(n1454), .C0(n1450), 
        .Y(n1451) );
  AOI31_X0P5M_A12TR U1567 ( .A0(n1454), .A1(n1453), .A2(n1452), .B0(n1451), 
        .Y(\outreg_stage2/N34 ) );
  ADDF_X1M_A12TR U1568 ( .A(in_s2[1]), .B(acc_s2[1]), .CI(n1455), .CO(n1456), 
        .S(out[1]) );
  ADDF_X1M_A12TR U1569 ( .A(in_s2[2]), .B(acc_s2[2]), .CI(n1456), .CO(n1457), 
        .S(out[2]) );
  ADDF_X1M_A12TR U1570 ( .A(in_s2[3]), .B(acc_s2[3]), .CI(n1457), .CO(n1458), 
        .S(out[3]) );
  ADDF_X1M_A12TR U1571 ( .A(in_s2[4]), .B(acc_s2[4]), .CI(n1458), .CO(n1459), 
        .S(out[4]) );
  ADDF_X1M_A12TR U1572 ( .A(in_s2[5]), .B(acc_s2[5]), .CI(n1459), .CO(n1460), 
        .S(out[5]) );
  ADDF_X1M_A12TR U1573 ( .A(in_s2[6]), .B(acc_s2[6]), .CI(n1460), .CO(n1461), 
        .S(out[6]) );
  ADDF_X1M_A12TR U1574 ( .A(in_s2[7]), .B(acc_s2[7]), .CI(n1461), .CO(n1462), 
        .S(out[7]) );
  ADDF_X1M_A12TR U1575 ( .A(in_s2[8]), .B(acc_s2[8]), .CI(n1462), .CO(n1463), 
        .S(out[8]) );
  ADDF_X1M_A12TR U1576 ( .A(in_s2[9]), .B(acc_s2[9]), .CI(n1463), .CO(n1464), 
        .S(out[9]) );
  ADDF_X1M_A12TR U1577 ( .A(in_s2[10]), .B(acc_s2[10]), .CI(n1464), .CO(n1465), 
        .S(out[10]) );
  ADDF_X1M_A12TR U1578 ( .A(in_s2[11]), .B(acc_s2[11]), .CI(n1465), .CO(n1466), 
        .S(out[11]) );
  ADDF_X1M_A12TR U1579 ( .A(in_s2[12]), .B(acc_s2[12]), .CI(n1466), .CO(n1467), 
        .S(out[12]) );
  ADDF_X1M_A12TR U1580 ( .A(in_s2[13]), .B(acc_s2[13]), .CI(n1467), .CO(n1468), 
        .S(out[13]) );
  ADDF_X1M_A12TR U1581 ( .A(in_s2[14]), .B(acc_s2[14]), .CI(n1468), .CO(n1469), 
        .S(out[14]) );
  ADDF_X1M_A12TR U1582 ( .A(in_s2[15]), .B(acc_s2[15]), .CI(n1469), .CO(n1470), 
        .S(out[15]) );
  ADDF_X1M_A12TR U1583 ( .A(in_s2[16]), .B(acc_s2[16]), .CI(n1470), .CO(n1471), 
        .S(out[16]) );
  ADDF_X1M_A12TR U1584 ( .A(in_s2[17]), .B(acc_s2[17]), .CI(n1471), .CO(n1472), 
        .S(out[17]) );
  ADDF_X1M_A12TR U1585 ( .A(in_s2[18]), .B(acc_s2[18]), .CI(n1472), .CO(n1473), 
        .S(out[18]) );
  ADDF_X1M_A12TR U1586 ( .A(in_s2[19]), .B(acc_s2[19]), .CI(n1473), .CO(n1474), 
        .S(out[19]) );
  ADDF_X1M_A12TR U1587 ( .A(in_s2[20]), .B(acc_s2[20]), .CI(n1474), .CO(n1475), 
        .S(out[20]) );
  ADDF_X1M_A12TR U1588 ( .A(in_s2[21]), .B(acc_s2[21]), .CI(n1475), .CO(n1476), 
        .S(out[21]) );
  ADDF_X1M_A12TR U1589 ( .A(in_s2[22]), .B(acc_s2[22]), .CI(n1476), .CO(n1477), 
        .S(out[22]) );
  ADDF_X1M_A12TR U1590 ( .A(in_s2[23]), .B(acc_s2[23]), .CI(n1477), .CO(n1478), 
        .S(out[23]) );
  ADDF_X1M_A12TR U1591 ( .A(in_s2[24]), .B(acc_s2[24]), .CI(n1478), .CO(n1479), 
        .S(out[24]) );
  ADDF_X1M_A12TR U1592 ( .A(in_s2[25]), .B(acc_s2[25]), .CI(n1479), .CO(n1480), 
        .S(out[25]) );
  ADDF_X1M_A12TR U1593 ( .A(in_s2[26]), .B(acc_s2[26]), .CI(n1480), .CO(n1481), 
        .S(out[26]) );
  ADDF_X1M_A12TR U1594 ( .A(in_s2[27]), .B(acc_s2[27]), .CI(n1481), .CO(n1482), 
        .S(out[27]) );
  ADDF_X1M_A12TR U1595 ( .A(in_s2[28]), .B(acc_s2[28]), .CI(n1482), .CO(n1483), 
        .S(out[28]) );
  ADDF_X1M_A12TR U1596 ( .A(in_s2[29]), .B(acc_s2[29]), .CI(n1483), .CO(n1484), 
        .S(out[29]) );
  ADDF_X1M_A12TR U1597 ( .A(in_s2[30]), .B(acc_s2[30]), .CI(n1484), .CO(n1272), 
        .S(out[30]) );
endmodule

`timescale 1ns / 1ps

module test;
  reg R1b, R2b;
  wire L2b, Ldb;
  reg trigger;
  reg nsR, npR;
  reg clk1;
  reg clk2;
  integer counter = 0;
 // wire clk1;
 // wire clk2;
  reg reset;
  reg [ 31 : 0 ] a;
  reg [ 31 : 0 ] b;
  wire [ 31 : 0 ] out;

  integer a_in[9:0];
  integer b_in[9:0];

  mul_add #( 32, 0 )dut (
    .clk1 ( clk1 ),
    .clk2 ( clk2 ),
    .reset ( reset ),
    .a ( a ),
    .b ( b ),
    .out ( out )
  );

  initial begin
     $sdf_annotate("Top.mapped.sdf", dut);
  end

  initial begin
     $prsim("afterclock.prs");

     $to_prsim ("nsR", "g._sReset");
     $to_prsim ("npR", "g._pReset");

     $from_prsim ( "L1.a", "clk1" );
     $from_prsim ( "L2.a", "clk2" );
     $from_prsim ( "L1.b", "trigger" );

  end
  initial begin

    counter = 0;
    a_in[0] = 10;
    a_in[1] = 3;
    a_in[2] = 10;
    a_in[3] = 2;
    a_in[4] = 15;
    a_in[5] = 100;
    a_in[6] = 39;
    a_in[7] = 101;
    a_in[8] = 22;
    a_in[9] = 151;

    b_in[0] = 7;
    b_in[1] = 10;
    b_in[2] = 1;
    b_in[3] = 12;
    b_in[4] = 10;
    b_in[5] = 7;
    b_in[6] = 10;
    b_in[7] = 1;
    b_in[8] = 12;
    b_in[9] = 10;

    nsR = 0;
    #90 npR = 1;
    #90 npR = 0;
    #90 npR = 1;
    #90 nsR <= 1;
    #30 reset = 1;
    #100 reset = 0;
    #1000 $finish;  
  end
 
  always @(posedge trigger) begin
          a = a_in[counter];
          b = b_in[counter]; 
  end
  
  always @(posedge clk1) begin
       if ( reset == 0 ) begin
          counter = counter + 1;
       end
  end 

  initial begin
    $dumpfile("mul_add.vcd");
    $dumpvars;
  end

  initial begin
    $display("\t\ttime,\treset,\tclk1,\tclk2,\t\ta,\t\tb,\t\ta_s1,\t\tb_s1,\t\tin_s2,\t\tacc_s2,\t\t\out");
    $monitor("%d,\t%b,\t%b,\t%d,\t%d,\t%d,\t%d,\t%d,\t%d,\t%d,\t%d",$time,reset,clk1,clk2,a,b,dut.a_s1,dut.b_s1,dut.in_s2,dut.acc_s2,out);
  end


endmodule 
